module image_rom_r (
    input  wire [4:0] row,
    input  wire [4:0] col,
    output reg [7:0] data
);

    reg [7:0] rom [0:31][0:31];

    initial begin
        rom[0][0] = 8'd167;
        rom[0][1] = 8'd167;
        rom[0][2] = 8'd169;
        rom[0][3] = 8'd173;
        rom[0][4] = 8'd177;
        rom[0][5] = 8'd180;
        rom[0][6] = 8'd182;
        rom[0][7] = 8'd185;
        rom[0][8] = 8'd187;
        rom[0][9] = 8'd189;
        rom[0][10] = 8'd192;
        rom[0][11] = 8'd196;
        rom[0][12] = 8'd200;
        rom[0][13] = 8'd204;
        rom[0][14] = 8'd207;
        rom[0][15] = 8'd210;
        rom[0][16] = 8'd212;
        rom[0][17] = 8'd212;
        rom[0][18] = 8'd213;
        rom[0][19] = 8'd214;
        rom[0][20] = 8'd217;
        rom[0][21] = 8'd221;
        rom[0][22] = 8'd225;
        rom[0][23] = 8'd226;
        rom[0][24] = 8'd226;
        rom[0][25] = 8'd228;
        rom[0][26] = 8'd230;
        rom[0][27] = 8'd232;
        rom[0][28] = 8'd232;
        rom[0][29] = 8'd233;
        rom[0][30] = 8'd235;
        rom[0][31] = 8'd234;
        rom[1][0] = 8'd171;
        rom[1][1] = 8'd171;
        rom[1][2] = 8'd173;
        rom[1][3] = 8'd176;
        rom[1][4] = 8'd179;
        rom[1][5] = 8'd182;
        rom[1][6] = 8'd185;
        rom[1][7] = 8'd189;
        rom[1][8] = 8'd191;
        rom[1][9] = 8'd193;
        rom[1][10] = 8'd196;
        rom[1][11] = 8'd199;
        rom[1][12] = 8'd203;
        rom[1][13] = 8'd207;
        rom[1][14] = 8'd210;
        rom[1][15] = 8'd213;
        rom[1][16] = 8'd215;
        rom[1][17] = 8'd216;
        rom[1][18] = 8'd215;
        rom[1][19] = 8'd217;
        rom[1][20] = 8'd218;
        rom[1][21] = 8'd228;
        rom[1][22] = 8'd233;
        rom[1][23] = 8'd227;
        rom[1][24] = 8'd228;
        rom[1][25] = 8'd229;
        rom[1][26] = 8'd231;
        rom[1][27] = 8'd233;
        rom[1][28] = 8'd232;
        rom[1][29] = 8'd233;
        rom[1][30] = 8'd234;
        rom[1][31] = 8'd233;
        rom[2][0] = 8'd175;
        rom[2][1] = 8'd175;
        rom[2][2] = 8'd178;
        rom[2][3] = 8'd181;
        rom[2][4] = 8'd183;
        rom[2][5] = 8'd187;
        rom[2][6] = 8'd190;
        rom[2][7] = 8'd194;
        rom[2][8] = 8'd195;
        rom[2][9] = 8'd197;
        rom[2][10] = 8'd200;
        rom[2][11] = 8'd204;
        rom[2][12] = 8'd208;
        rom[2][13] = 8'd212;
        rom[2][14] = 8'd215;
        rom[2][15] = 8'd217;
        rom[2][16] = 8'd219;
        rom[2][17] = 8'd221;
        rom[2][18] = 8'd220;
        rom[2][19] = 8'd220;
        rom[2][20] = 8'd223;
        rom[2][21] = 8'd230;
        rom[2][22] = 8'd234;
        rom[2][23] = 8'd231;
        rom[2][24] = 8'd231;
        rom[2][25] = 8'd232;
        rom[2][26] = 8'd235;
        rom[2][27] = 8'd236;
        rom[2][28] = 8'd235;
        rom[2][29] = 8'd235;
        rom[2][30] = 8'd235;
        rom[2][31] = 8'd234;
        rom[3][0] = 8'd179;
        rom[3][1] = 8'd179;
        rom[3][2] = 8'd183;
        rom[3][3] = 8'd187;
        rom[3][4] = 8'd189;
        rom[3][5] = 8'd192;
        rom[3][6] = 8'd196;
        rom[3][7] = 8'd199;
        rom[3][8] = 8'd200;
        rom[3][9] = 8'd201;
        rom[3][10] = 8'd204;
        rom[3][11] = 8'd207;
        rom[3][12] = 8'd211;
        rom[3][13] = 8'd216;
        rom[3][14] = 8'd219;
        rom[3][15] = 8'd221;
        rom[3][16] = 8'd222;
        rom[3][17] = 8'd223;
        rom[3][18] = 8'd223;
        rom[3][19] = 8'd224;
        rom[3][20] = 8'd226;
        rom[3][21] = 8'd228;
        rom[3][22] = 8'd230;
        rom[3][23] = 8'd233;
        rom[3][24] = 8'd234;
        rom[3][25] = 8'd235;
        rom[3][26] = 8'd238;
        rom[3][27] = 8'd240;
        rom[3][28] = 8'd237;
        rom[3][29] = 8'd236;
        rom[3][30] = 8'd235;
        rom[3][31] = 8'd235;
        rom[4][0] = 8'd183;
        rom[4][1] = 8'd184;
        rom[4][2] = 8'd187;
        rom[4][3] = 8'd191;
        rom[4][4] = 8'd193;
        rom[4][5] = 8'd196;
        rom[4][6] = 8'd200;
        rom[4][7] = 8'd203;
        rom[4][8] = 8'd204;
        rom[4][9] = 8'd205;
        rom[4][10] = 8'd207;
        rom[4][11] = 8'd211;
        rom[4][12] = 8'd215;
        rom[4][13] = 8'd220;
        rom[4][14] = 8'd222;
        rom[4][15] = 8'd224;
        rom[4][16] = 8'd225;
        rom[4][17] = 8'd226;
        rom[4][18] = 8'd227;
        rom[4][19] = 8'd228;
        rom[4][20] = 8'd229;
        rom[4][21] = 8'd232;
        rom[4][22] = 8'd233;
        rom[4][23] = 8'd234;
        rom[4][24] = 8'd235;
        rom[4][25] = 8'd235;
        rom[4][26] = 8'd239;
        rom[4][27] = 8'd240;
        rom[4][28] = 8'd238;
        rom[4][29] = 8'd237;
        rom[4][30] = 8'd235;
        rom[4][31] = 8'd235;
        rom[5][0] = 8'd188;
        rom[5][1] = 8'd189;
        rom[5][2] = 8'd193;
        rom[5][3] = 8'd196;
        rom[5][4] = 8'd198;
        rom[5][5] = 8'd201;
        rom[5][6] = 8'd204;
        rom[5][7] = 8'd207;
        rom[5][8] = 8'd207;
        rom[5][9] = 8'd208;
        rom[5][10] = 8'd210;
        rom[5][11] = 8'd214;
        rom[5][12] = 8'd218;
        rom[5][13] = 8'd223;
        rom[5][14] = 8'd224;
        rom[5][15] = 8'd226;
        rom[5][16] = 8'd226;
        rom[5][17] = 8'd227;
        rom[5][18] = 8'd230;
        rom[5][19] = 8'd232;
        rom[5][20] = 8'd234;
        rom[5][21] = 8'd236;
        rom[5][22] = 8'd236;
        rom[5][23] = 8'd236;
        rom[5][24] = 8'd236;
        rom[5][25] = 8'd236;
        rom[5][26] = 8'd238;
        rom[5][27] = 8'd238;
        rom[5][28] = 8'd238;
        rom[5][29] = 8'd237;
        rom[5][30] = 8'd236;
        rom[5][31] = 8'd236;
        rom[6][0] = 8'd194;
        rom[6][1] = 8'd195;
        rom[6][2] = 8'd199;
        rom[6][3] = 8'd202;
        rom[6][4] = 8'd204;
        rom[6][5] = 8'd206;
        rom[6][6] = 8'd208;
        rom[6][7] = 8'd210;
        rom[6][8] = 8'd211;
        rom[6][9] = 8'd215;
        rom[6][10] = 8'd218;
        rom[6][11] = 8'd222;
        rom[6][12] = 8'd227;
        rom[6][13] = 8'd232;
        rom[6][14] = 8'd233;
        rom[6][15] = 8'd234;
        rom[6][16] = 8'd236;
        rom[6][17] = 8'd238;
        rom[6][18] = 8'd240;
        rom[6][19] = 8'd239;
        rom[6][20] = 8'd239;
        rom[6][21] = 8'd240;
        rom[6][22] = 8'd239;
        rom[6][23] = 8'd238;
        rom[6][24] = 8'd238;
        rom[6][25] = 8'd238;
        rom[6][26] = 8'd239;
        rom[6][27] = 8'd240;
        rom[6][28] = 8'd240;
        rom[6][29] = 8'd239;
        rom[6][30] = 8'd238;
        rom[6][31] = 8'd238;
        rom[7][0] = 8'd200;
        rom[7][1] = 8'd202;
        rom[7][2] = 8'd205;
        rom[7][3] = 8'd209;
        rom[7][4] = 8'd210;
        rom[7][5] = 8'd212;
        rom[7][6] = 8'd213;
        rom[7][7] = 8'd213;
        rom[7][8] = 8'd216;
        rom[7][9] = 8'd212;
        rom[7][10] = 8'd208;
        rom[7][11] = 8'd209;
        rom[7][12] = 8'd210;
        rom[7][13] = 8'd210;
        rom[7][14] = 8'd212;
        rom[7][15] = 8'd213;
        rom[7][16] = 8'd213;
        rom[7][17] = 8'd213;
        rom[7][18] = 8'd222;
        rom[7][19] = 8'd242;
        rom[7][20] = 8'd243;
        rom[7][21] = 8'd236;
        rom[7][22] = 8'd238;
        rom[7][23] = 8'd242;
        rom[7][24] = 8'd241;
        rom[7][25] = 8'd241;
        rom[7][26] = 8'd242;
        rom[7][27] = 8'd242;
        rom[7][28] = 8'd242;
        rom[7][29] = 8'd242;
        rom[7][30] = 8'd241;
        rom[7][31] = 8'd241;
        rom[8][0] = 8'd204;
        rom[8][1] = 8'd208;
        rom[8][2] = 8'd212;
        rom[8][3] = 8'd215;
        rom[8][4] = 8'd216;
        rom[8][5] = 8'd217;
        rom[8][6] = 8'd218;
        rom[8][7] = 8'd220;
        rom[8][8] = 8'd222;
        rom[8][9] = 8'd152;
        rom[8][10] = 8'd118;
        rom[8][11] = 8'd120;
        rom[8][12] = 8'd116;
        rom[8][13] = 8'd117;
        rom[8][14] = 8'd120;
        rom[8][15] = 8'd126;
        rom[8][16] = 8'd132;
        rom[8][17] = 8'd133;
        rom[8][18] = 8'd154;
        rom[8][19] = 8'd207;
        rom[8][20] = 8'd212;
        rom[8][21] = 8'd203;
        rom[8][22] = 8'd230;
        rom[8][23] = 8'd247;
        rom[8][24] = 8'd244;
        rom[8][25] = 8'd244;
        rom[8][26] = 8'd244;
        rom[8][27] = 8'd245;
        rom[8][28] = 8'd245;
        rom[8][29] = 8'd244;
        rom[8][30] = 8'd243;
        rom[8][31] = 8'd243;
        rom[9][0] = 8'd205;
        rom[9][1] = 8'd199;
        rom[9][2] = 8'd216;
        rom[9][3] = 8'd221;
        rom[9][4] = 8'd222;
        rom[9][5] = 8'd222;
        rom[9][6] = 8'd223;
        rom[9][7] = 8'd226;
        rom[9][8] = 8'd225;
        rom[9][9] = 8'd128;
        rom[9][10] = 8'd96;
        rom[9][11] = 8'd101;
        rom[9][12] = 8'd102;
        rom[9][13] = 8'd103;
        rom[9][14] = 8'd104;
        rom[9][15] = 8'd110;
        rom[9][16] = 8'd121;
        rom[9][17] = 8'd125;
        rom[9][18] = 8'd149;
        rom[9][19] = 8'd183;
        rom[9][20] = 8'd186;
        rom[9][21] = 8'd193;
        rom[9][22] = 8'd219;
        rom[9][23] = 8'd232;
        rom[9][24] = 8'd234;
        rom[9][25] = 8'd244;
        rom[9][26] = 8'd247;
        rom[9][27] = 8'd247;
        rom[9][28] = 8'd247;
        rom[9][29] = 8'd247;
        rom[9][30] = 8'd246;
        rom[9][31] = 8'd247;
        rom[10][0] = 8'd188;
        rom[10][1] = 8'd192;
        rom[10][2] = 8'd223;
        rom[10][3] = 8'd225;
        rom[10][4] = 8'd228;
        rom[10][5] = 8'd228;
        rom[10][6] = 8'd228;
        rom[10][7] = 8'd231;
        rom[10][8] = 8'd225;
        rom[10][9] = 8'd132;
        rom[10][10] = 8'd103;
        rom[10][11] = 8'd107;
        rom[10][12] = 8'd107;
        rom[10][13] = 8'd105;
        rom[10][14] = 8'd110;
        rom[10][15] = 8'd117;
        rom[10][16] = 8'd125;
        rom[10][17] = 8'd131;
        rom[10][18] = 8'd145;
        rom[10][19] = 8'd186;
        rom[10][20] = 8'd183;
        rom[10][21] = 8'd152;
        rom[10][22] = 8'd168;
        rom[10][23] = 8'd169;
        rom[10][24] = 8'd176;
        rom[10][25] = 8'd224;
        rom[10][26] = 8'd249;
        rom[10][27] = 8'd251;
        rom[10][28] = 8'd251;
        rom[10][29] = 8'd251;
        rom[10][30] = 8'd249;
        rom[10][31] = 8'd248;
        rom[11][0] = 8'd105;
        rom[11][1] = 8'd163;
        rom[11][2] = 8'd201;
        rom[11][3] = 8'd229;
        rom[11][4] = 8'd233;
        rom[11][5] = 8'd235;
        rom[11][6] = 8'd235;
        rom[11][7] = 8'd237;
        rom[11][8] = 8'd229;
        rom[11][9] = 8'd139;
        rom[11][10] = 8'd107;
        rom[11][11] = 8'd108;
        rom[11][12] = 8'd98;
        rom[11][13] = 8'd96;
        rom[11][14] = 8'd107;
        rom[11][15] = 8'd118;
        rom[11][16] = 8'd129;
        rom[11][17] = 8'd133;
        rom[11][18] = 8'd140;
        rom[11][19] = 8'd178;
        rom[11][20] = 8'd169;
        rom[11][21] = 8'd121;
        rom[11][22] = 8'd117;
        rom[11][23] = 8'd134;
        rom[11][24] = 8'd144;
        rom[11][25] = 8'd174;
        rom[11][26] = 8'd239;
        rom[11][27] = 8'd245;
        rom[11][28] = 8'd242;
        rom[11][29] = 8'd241;
        rom[11][30] = 8'd242;
        rom[11][31] = 8'd227;
        rom[12][0] = 8'd61;
        rom[12][1] = 8'd97;
        rom[12][2] = 8'd109;
        rom[12][3] = 8'd203;
        rom[12][4] = 8'd241;
        rom[12][5] = 8'd239;
        rom[12][6] = 8'd240;
        rom[12][7] = 8'd238;
        rom[12][8] = 8'd233;
        rom[12][9] = 8'd148;
        rom[12][10] = 8'd116;
        rom[12][11] = 8'd113;
        rom[12][12] = 8'd96;
        rom[12][13] = 8'd97;
        rom[12][14] = 8'd108;
        rom[12][15] = 8'd119;
        rom[12][16] = 8'd132;
        rom[12][17] = 8'd142;
        rom[12][18] = 8'd153;
        rom[12][19] = 8'd180;
        rom[12][20] = 8'd165;
        rom[12][21] = 8'd120;
        rom[12][22] = 8'd132;
        rom[12][23] = 8'd143;
        rom[12][24] = 8'd139;
        rom[12][25] = 8'd150;
        rom[12][26] = 8'd224;
        rom[12][27] = 8'd193;
        rom[12][28] = 8'd199;
        rom[12][29] = 8'd191;
        rom[12][30] = 8'd199;
        rom[12][31] = 8'd180;
        rom[13][0] = 8'd56;
        rom[13][1] = 8'd67;
        rom[13][2] = 8'd61;
        rom[13][3] = 8'd172;
        rom[13][4] = 8'd248;
        rom[13][5] = 8'd248;
        rom[13][6] = 8'd249;
        rom[13][7] = 8'd168;
        rom[13][8] = 8'd197;
        rom[13][9] = 8'd138;
        rom[13][10] = 8'd116;
        rom[13][11] = 8'd113;
        rom[13][12] = 8'd96;
        rom[13][13] = 8'd99;
        rom[13][14] = 8'd108;
        rom[13][15] = 8'd119;
        rom[13][16] = 8'd133;
        rom[13][17] = 8'd136;
        rom[13][18] = 8'd148;
        rom[13][19] = 8'd174;
        rom[13][20] = 8'd160;
        rom[13][21] = 8'd123;
        rom[13][22] = 8'd170;
        rom[13][23] = 8'd153;
        rom[13][24] = 8'd115;
        rom[13][25] = 8'd141;
        rom[13][26] = 8'd180;
        rom[13][27] = 8'd127;
        rom[13][28] = 8'd128;
        rom[13][29] = 8'd129;
        rom[13][30] = 8'd144;
        rom[13][31] = 8'd135;
        rom[14][0] = 8'd88;
        rom[14][1] = 8'd90;
        rom[14][2] = 8'd90;
        rom[14][3] = 8'd132;
        rom[14][4] = 8'd176;
        rom[14][5] = 8'd188;
        rom[14][6] = 8'd188;
        rom[14][7] = 8'd120;
        rom[14][8] = 8'd139;
        rom[14][9] = 8'd122;
        rom[14][10] = 8'd122;
        rom[14][11] = 8'd111;
        rom[14][12] = 8'd92;
        rom[14][13] = 8'd93;
        rom[14][14] = 8'd104;
        rom[14][15] = 8'd114;
        rom[14][16] = 8'd129;
        rom[14][17] = 8'd129;
        rom[14][18] = 8'd129;
        rom[14][19] = 8'd159;
        rom[14][20] = 8'd160;
        rom[14][21] = 8'd153;
        rom[14][22] = 8'd192;
        rom[14][23] = 8'd179;
        rom[14][24] = 8'd126;
        rom[14][25] = 8'd128;
        rom[14][26] = 8'd154;
        rom[14][27] = 8'd115;
        rom[14][28] = 8'd123;
        rom[14][29] = 8'd130;
        rom[14][30] = 8'd163;
        rom[14][31] = 8'd165;
        rom[15][0] = 8'd126;
        rom[15][1] = 8'd124;
        rom[15][2] = 8'd131;
        rom[15][3] = 8'd125;
        rom[15][4] = 8'd126;
        rom[15][5] = 8'd133;
        rom[15][6] = 8'd137;
        rom[15][7] = 8'd142;
        rom[15][8] = 8'd138;
        rom[15][9] = 8'd112;
        rom[15][10] = 8'd116;
        rom[15][11] = 8'd103;
        rom[15][12] = 8'd91;
        rom[15][13] = 8'd90;
        rom[15][14] = 8'd99;
        rom[15][15] = 8'd109;
        rom[15][16] = 8'd118;
        rom[15][17] = 8'd129;
        rom[15][18] = 8'd127;
        rom[15][19] = 8'd161;
        rom[15][20] = 8'd194;
        rom[15][21] = 8'd179;
        rom[15][22] = 8'd187;
        rom[15][23] = 8'd189;
        rom[15][24] = 8'd136;
        rom[15][25] = 8'd156;
        rom[15][26] = 8'd172;
        rom[15][27] = 8'd197;
        rom[15][28] = 8'd205;
        rom[15][29] = 8'd203;
        rom[15][30] = 8'd208;
        rom[15][31] = 8'd195;
        rom[16][0] = 8'd150;
        rom[16][1] = 8'd160;
        rom[16][2] = 8'd164;
        rom[16][3] = 8'd167;
        rom[16][4] = 8'd171;
        rom[16][5] = 8'd174;
        rom[16][6] = 8'd177;
        rom[16][7] = 8'd181;
        rom[16][8] = 8'd172;
        rom[16][9] = 8'd110;
        rom[16][10] = 8'd95;
        rom[16][11] = 8'd94;
        rom[16][12] = 8'd91;
        rom[16][13] = 8'd91;
        rom[16][14] = 8'd99;
        rom[16][15] = 8'd105;
        rom[16][16] = 8'd108;
        rom[16][17] = 8'd118;
        rom[16][18] = 8'd125;
        rom[16][19] = 8'd182;
        rom[16][20] = 8'd197;
        rom[16][21] = 8'd177;
        rom[16][22] = 8'd196;
        rom[16][23] = 8'd161;
        rom[16][24] = 8'd138;
        rom[16][25] = 8'd163;
        rom[16][26] = 8'd170;
        rom[16][27] = 8'd240;
        rom[16][28] = 8'd232;
        rom[16][29] = 8'd213;
        rom[16][30] = 8'd182;
        rom[16][31] = 8'd184;
        rom[17][0] = 8'd156;
        rom[17][1] = 8'd162;
        rom[17][2] = 8'd163;
        rom[17][3] = 8'd165;
        rom[17][4] = 8'd166;
        rom[17][5] = 8'd170;
        rom[17][6] = 8'd174;
        rom[17][7] = 8'd180;
        rom[17][8] = 8'd168;
        rom[17][9] = 8'd105;
        rom[17][10] = 8'd89;
        rom[17][11] = 8'd91;
        rom[17][12] = 8'd93;
        rom[17][13] = 8'd93;
        rom[17][14] = 8'd100;
        rom[17][15] = 8'd106;
        rom[17][16] = 8'd104;
        rom[17][17] = 8'd111;
        rom[17][18] = 8'd120;
        rom[17][19] = 8'd170;
        rom[17][20] = 8'd168;
        rom[17][21] = 8'd199;
        rom[17][22] = 8'd176;
        rom[17][23] = 8'd133;
        rom[17][24] = 8'd119;
        rom[17][25] = 8'd112;
        rom[17][26] = 8'd154;
        rom[17][27] = 8'd218;
        rom[17][28] = 8'd215;
        rom[17][29] = 8'd183;
        rom[17][30] = 8'd167;
        rom[17][31] = 8'd175;
        rom[18][0] = 8'd152;
        rom[18][1] = 8'd154;
        rom[18][2] = 8'd158;
        rom[18][3] = 8'd164;
        rom[18][4] = 8'd167;
        rom[18][5] = 8'd168;
        rom[18][6] = 8'd169;
        rom[18][7] = 8'd171;
        rom[18][8] = 8'd157;
        rom[18][9] = 8'd101;
        rom[18][10] = 8'd86;
        rom[18][11] = 8'd84;
        rom[18][12] = 8'd101;
        rom[18][13] = 8'd114;
        rom[18][14] = 8'd104;
        rom[18][15] = 8'd100;
        rom[18][16] = 8'd101;
        rom[18][17] = 8'd108;
        rom[18][18] = 8'd117;
        rom[18][19] = 8'd150;
        rom[18][20] = 8'd197;
        rom[18][21] = 8'd191;
        rom[18][22] = 8'd143;
        rom[18][23] = 8'd111;
        rom[18][24] = 8'd89;
        rom[18][25] = 8'd86;
        rom[18][26] = 8'd145;
        rom[18][27] = 8'd210;
        rom[18][28] = 8'd203;
        rom[18][29] = 8'd166;
        rom[18][30] = 8'd164;
        rom[18][31] = 8'd164;
        rom[19][0] = 8'd153;
        rom[19][1] = 8'd153;
        rom[19][2] = 8'd151;
        rom[19][3] = 8'd150;
        rom[19][4] = 8'd151;
        rom[19][5] = 8'd152;
        rom[19][6] = 8'd156;
        rom[19][7] = 8'd161;
        rom[19][8] = 8'd154;
        rom[19][9] = 8'd97;
        rom[19][10] = 8'd85;
        rom[19][11] = 8'd84;
        rom[19][12] = 8'd104;
        rom[19][13] = 8'd123;
        rom[19][14] = 8'd105;
        rom[19][15] = 8'd92;
        rom[19][16] = 8'd96;
        rom[19][17] = 8'd100;
        rom[19][18] = 8'd119;
        rom[19][19] = 8'd146;
        rom[19][20] = 8'd163;
        rom[19][21] = 8'd132;
        rom[19][22] = 8'd125;
        rom[19][23] = 8'd126;
        rom[19][24] = 8'd84;
        rom[19][25] = 8'd91;
        rom[19][26] = 8'd167;
        rom[19][27] = 8'd208;
        rom[19][28] = 8'd182;
        rom[19][29] = 8'd152;
        rom[19][30] = 8'd160;
        rom[19][31] = 8'd156;
        rom[20][0] = 8'd138;
        rom[20][1] = 8'd139;
        rom[20][2] = 8'd145;
        rom[20][3] = 8'd151;
        rom[20][4] = 8'd155;
        rom[20][5] = 8'd162;
        rom[20][6] = 8'd170;
        rom[20][7] = 8'd174;
        rom[20][8] = 8'd163;
        rom[20][9] = 8'd94;
        rom[20][10] = 8'd87;
        rom[20][11] = 8'd84;
        rom[20][12] = 8'd92;
        rom[20][13] = 8'd110;
        rom[20][14] = 8'd96;
        rom[20][15] = 8'd84;
        rom[20][16] = 8'd92;
        rom[20][17] = 8'd96;
        rom[20][18] = 8'd112;
        rom[20][19] = 8'd128;
        rom[20][20] = 8'd116;
        rom[20][21] = 8'd89;
        rom[20][22] = 8'd126;
        rom[20][23] = 8'd111;
        rom[20][24] = 8'd75;
        rom[20][25] = 8'd123;
        rom[20][26] = 8'd201;
        rom[20][27] = 8'd203;
        rom[20][28] = 8'd160;
        rom[20][29] = 8'd142;
        rom[20][30] = 8'd153;
        rom[20][31] = 8'd152;
        rom[21][0] = 8'd152;
        rom[21][1] = 8'd158;
        rom[21][2] = 8'd160;
        rom[21][3] = 8'd165;
        rom[21][4] = 8'd165;
        rom[21][5] = 8'd161;
        rom[21][6] = 8'd160;
        rom[21][7] = 8'd161;
        rom[21][8] = 8'd153;
        rom[21][9] = 8'd98;
        rom[21][10] = 8'd76;
        rom[21][11] = 8'd73;
        rom[21][12] = 8'd74;
        rom[21][13] = 8'd82;
        rom[21][14] = 8'd81;
        rom[21][15] = 8'd80;
        rom[21][16] = 8'd89;
        rom[21][17] = 8'd92;
        rom[21][18] = 8'd94;
        rom[21][19] = 8'd112;
        rom[21][20] = 8'd111;
        rom[21][21] = 8'd88;
        rom[21][22] = 8'd129;
        rom[21][23] = 8'd107;
        rom[21][24] = 8'd116;
        rom[21][25] = 8'd174;
        rom[21][26] = 8'd206;
        rom[21][27] = 8'd188;
        rom[21][28] = 8'd149;
        rom[21][29] = 8'd155;
        rom[21][30] = 8'd155;
        rom[21][31] = 8'd151;
        rom[22][0] = 8'd152;
        rom[22][1] = 8'd151;
        rom[22][2] = 8'd150;
        rom[22][3] = 8'd149;
        rom[22][4] = 8'd146;
        rom[22][5] = 8'd145;
        rom[22][6] = 8'd148;
        rom[22][7] = 8'd151;
        rom[22][8] = 8'd145;
        rom[22][9] = 8'd89;
        rom[22][10] = 8'd65;
        rom[22][11] = 8'd65;
        rom[22][12] = 8'd54;
        rom[22][13] = 8'd58;
        rom[22][14] = 8'd64;
        rom[22][15] = 8'd65;
        rom[22][16] = 8'd71;
        rom[22][17] = 8'd77;
        rom[22][18] = 8'd85;
        rom[22][19] = 8'd106;
        rom[22][20] = 8'd88;
        rom[22][21] = 8'd87;
        rom[22][22] = 8'd117;
        rom[22][23] = 8'd149;
        rom[22][24] = 8'd190;
        rom[22][25] = 8'd202;
        rom[22][26] = 8'd200;
        rom[22][27] = 8'd168;
        rom[22][28] = 8'd140;
        rom[22][29] = 8'd154;
        rom[22][30] = 8'd157;
        rom[22][31] = 8'd152;
        rom[23][0] = 8'd135;
        rom[23][1] = 8'd130;
        rom[23][2] = 8'd132;
        rom[23][3] = 8'd133;
        rom[23][4] = 8'd138;
        rom[23][5] = 8'd142;
        rom[23][6] = 8'd147;
        rom[23][7] = 8'd145;
        rom[23][8] = 8'd118;
        rom[23][9] = 8'd68;
        rom[23][10] = 8'd64;
        rom[23][11] = 8'd64;
        rom[23][12] = 8'd48;
        rom[23][13] = 8'd69;
        rom[23][14] = 8'd69;
        rom[23][15] = 8'd66;
        rom[23][16] = 8'd71;
        rom[23][17] = 8'd68;
        rom[23][18] = 8'd79;
        rom[23][19] = 8'd104;
        rom[23][20] = 8'd74;
        rom[23][21] = 8'd71;
        rom[23][22] = 8'd113;
        rom[23][23] = 8'd189;
        rom[23][24] = 8'd207;
        rom[23][25] = 8'd204;
        rom[23][26] = 8'd190;
        rom[23][27] = 8'd153;
        rom[23][28] = 8'd144;
        rom[23][29] = 8'd152;
        rom[23][30] = 8'd157;
        rom[23][31] = 8'd149;
        rom[24][0] = 8'd132;
        rom[24][1] = 8'd128;
        rom[24][2] = 8'd129;
        rom[24][3] = 8'd128;
        rom[24][4] = 8'd136;
        rom[24][5] = 8'd142;
        rom[24][6] = 8'd144;
        rom[24][7] = 8'd125;
        rom[24][8] = 8'd102;
        rom[24][9] = 8'd87;
        rom[24][10] = 8'd68;
        rom[24][11] = 8'd47;
        rom[24][12] = 8'd35;
        rom[24][13] = 8'd62;
        rom[24][14] = 8'd60;
        rom[24][15] = 8'd52;
        rom[24][16] = 8'd64;
        rom[24][17] = 8'd69;
        rom[24][18] = 8'd68;
        rom[24][19] = 8'd72;
        rom[24][20] = 8'd49;
        rom[24][21] = 8'd84;
        rom[24][22] = 8'd177;
        rom[24][23] = 8'd207;
        rom[24][24] = 8'd202;
        rom[24][25] = 8'd199;
        rom[24][26] = 8'd170;
        rom[24][27] = 8'd134;
        rom[24][28] = 8'd147;
        rom[24][29] = 8'd151;
        rom[24][30] = 8'd161;
        rom[24][31] = 8'd147;
        rom[25][0] = 8'd128;
        rom[25][1] = 8'd128;
        rom[25][2] = 8'd133;
        rom[25][3] = 8'd132;
        rom[25][4] = 8'd135;
        rom[25][5] = 8'd140;
        rom[25][6] = 8'd136;
        rom[25][7] = 8'd124;
        rom[25][8] = 8'd107;
        rom[25][9] = 8'd71;
        rom[25][10] = 8'd48;
        rom[25][11] = 8'd36;
        rom[25][12] = 8'd26;
        rom[25][13] = 8'd27;
        rom[25][14] = 8'd29;
        rom[25][15] = 8'd29;
        rom[25][16] = 8'd30;
        rom[25][17] = 8'd41;
        rom[25][18] = 8'd38;
        rom[25][19] = 8'd35;
        rom[25][20] = 8'd49;
        rom[25][21] = 8'd146;
        rom[25][22] = 8'd200;
        rom[25][23] = 8'd199;
        rom[25][24] = 8'd199;
        rom[25][25] = 8'd192;
        rom[25][26] = 8'd145;
        rom[25][27] = 8'd137;
        rom[25][28] = 8'd148;
        rom[25][29] = 8'd153;
        rom[25][30] = 8'd158;
        rom[25][31] = 8'd148;
        rom[26][0] = 8'd126;
        rom[26][1] = 8'd128;
        rom[26][2] = 8'd132;
        rom[26][3] = 8'd135;
        rom[26][4] = 8'd131;
        rom[26][5] = 8'd116;
        rom[26][6] = 8'd95;
        rom[26][7] = 8'd71;
        rom[26][8] = 8'd52;
        rom[26][9] = 8'd37;
        rom[26][10] = 8'd37;
        rom[26][11] = 8'd35;
        rom[26][12] = 8'd30;
        rom[26][13] = 8'd31;
        rom[26][14] = 8'd27;
        rom[26][15] = 8'd28;
        rom[26][16] = 8'd27;
        rom[26][17] = 8'd33;
        rom[26][18] = 8'd39;
        rom[26][19] = 8'd57;
        rom[26][20] = 8'd130;
        rom[26][21] = 8'd190;
        rom[26][22] = 8'd190;
        rom[26][23] = 8'd195;
        rom[26][24] = 8'd198;
        rom[26][25] = 8'd176;
        rom[26][26] = 8'd124;
        rom[26][27] = 8'd111;
        rom[26][28] = 8'd122;
        rom[26][29] = 8'd155;
        rom[26][30] = 8'd153;
        rom[26][31] = 8'd145;
        rom[27][0] = 8'd126;
        rom[27][1] = 8'd127;
        rom[27][2] = 8'd127;
        rom[27][3] = 8'd114;
        rom[27][4] = 8'd91;
        rom[27][5] = 8'd66;
        rom[27][6] = 8'd46;
        rom[27][7] = 8'd41;
        rom[27][8] = 8'd42;
        rom[27][9] = 8'd39;
        rom[27][10] = 8'd35;
        rom[27][11] = 8'd34;
        rom[27][12] = 8'd35;
        rom[27][13] = 8'd45;
        rom[27][14] = 8'd37;
        rom[27][15] = 8'd31;
        rom[27][16] = 8'd34;
        rom[27][17] = 8'd35;
        rom[27][18] = 8'd58;
        rom[27][19] = 8'd130;
        rom[27][20] = 8'd174;
        rom[27][21] = 8'd186;
        rom[27][22] = 8'd188;
        rom[27][23] = 8'd191;
        rom[27][24] = 8'd190;
        rom[27][25] = 8'd148;
        rom[27][26] = 8'd119;
        rom[27][27] = 8'd122;
        rom[27][28] = 8'd120;
        rom[27][29] = 8'd146;
        rom[27][30] = 8'd147;
        rom[27][31] = 8'd137;
        rom[28][0] = 8'd121;
        rom[28][1] = 8'd113;
        rom[28][2] = 8'd90;
        rom[28][3] = 8'd64;
        rom[28][4] = 8'd46;
        rom[28][5] = 8'd41;
        rom[28][6] = 8'd40;
        rom[28][7] = 8'd41;
        rom[28][8] = 8'd40;
        rom[28][9] = 8'd38;
        rom[28][10] = 8'd33;
        rom[28][11] = 8'd31;
        rom[28][12] = 8'd34;
        rom[28][13] = 8'd44;
        rom[28][14] = 8'd41;
        rom[28][15] = 8'd37;
        rom[28][16] = 8'd41;
        rom[28][17] = 8'd46;
        rom[28][18] = 8'd114;
        rom[28][19] = 8'd176;
        rom[28][20] = 8'd175;
        rom[28][21] = 8'd181;
        rom[28][22] = 8'd187;
        rom[28][23] = 8'd188;
        rom[28][24] = 8'd174;
        rom[28][25] = 8'd121;
        rom[28][26] = 8'd115;
        rom[28][27] = 8'd139;
        rom[28][28] = 8'd158;
        rom[28][29] = 8'd150;
        rom[28][30] = 8'd140;
        rom[28][31] = 8'd134;
        rom[29][0] = 8'd88;
        rom[29][1] = 8'd65;
        rom[29][2] = 8'd46;
        rom[29][3] = 8'd42;
        rom[29][4] = 8'd40;
        rom[29][5] = 8'd39;
        rom[29][6] = 8'd40;
        rom[29][7] = 8'd39;
        rom[29][8] = 8'd39;
        rom[29][9] = 8'd39;
        rom[29][10] = 8'd36;
        rom[29][11] = 8'd33;
        rom[29][12] = 8'd34;
        rom[29][13] = 8'd39;
        rom[29][14] = 8'd37;
        rom[29][15] = 8'd38;
        rom[29][16] = 8'd64;
        rom[29][17] = 8'd124;
        rom[29][18] = 8'd167;
        rom[29][19] = 8'd178;
        rom[29][20] = 8'd178;
        rom[29][21] = 8'd182;
        rom[29][22] = 8'd185;
        rom[29][23] = 8'd184;
        rom[29][24] = 8'd152;
        rom[29][25] = 8'd114;
        rom[29][26] = 8'd120;
        rom[29][27] = 8'd143;
        rom[29][28] = 8'd150;
        rom[29][29] = 8'd138;
        rom[29][30] = 8'd127;
        rom[29][31] = 8'd125;
        rom[30][0] = 8'd44;
        rom[30][1] = 8'd36;
        rom[30][2] = 8'd36;
        rom[30][3] = 8'd41;
        rom[30][4] = 8'd39;
        rom[30][5] = 8'd35;
        rom[30][6] = 8'd37;
        rom[30][7] = 8'd40;
        rom[30][8] = 8'd40;
        rom[30][9] = 8'd39;
        rom[30][10] = 8'd37;
        rom[30][11] = 8'd38;
        rom[30][12] = 8'd40;
        rom[30][13] = 8'd39;
        rom[30][14] = 8'd37;
        rom[30][15] = 8'd62;
        rom[30][16] = 8'd134;
        rom[30][17] = 8'd181;
        rom[30][18] = 8'd182;
        rom[30][19] = 8'd177;
        rom[30][20] = 8'd177;
        rom[30][21] = 8'd181;
        rom[30][22] = 8'd180;
        rom[30][23] = 8'd169;
        rom[30][24] = 8'd121;
        rom[30][25] = 8'd127;
        rom[30][26] = 8'd131;
        rom[30][27] = 8'd139;
        rom[30][28] = 8'd147;
        rom[30][29] = 8'd132;
        rom[30][30] = 8'd120;
        rom[30][31] = 8'd124;
        rom[31][0] = 8'd39;
        rom[31][1] = 8'd36;
        rom[31][2] = 8'd37;
        rom[31][3] = 8'd41;
        rom[31][4] = 8'd39;
        rom[31][5] = 8'd35;
        rom[31][6] = 8'd37;
        rom[31][7] = 8'd41;
        rom[31][8] = 8'd42;
        rom[31][9] = 8'd40;
        rom[31][10] = 8'd38;
        rom[31][11] = 8'd41;
        rom[31][12] = 8'd43;
        rom[31][13] = 8'd50;
        rom[31][14] = 8'd91;
        rom[31][15] = 8'd141;
        rom[31][16] = 8'd167;
        rom[31][17] = 8'd177;
        rom[31][18] = 8'd181;
        rom[31][19] = 8'd175;
        rom[31][20] = 8'd178;
        rom[31][21] = 8'd176;
        rom[31][22] = 8'd174;
        rom[31][23] = 8'd143;
        rom[31][24] = 8'd117;
        rom[31][25] = 8'd140;
        rom[31][26] = 8'd133;
        rom[31][27] = 8'd109;
        rom[31][28] = 8'd115;
        rom[31][29] = 8'd116;
        rom[31][30] = 8'd120;
        rom[31][31] = 8'd128;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
