`timescale 1ns / 1ps

module conv2d_q17_top #(
    parameter WIDTH    = 32,
    parameter HEIGHT   = 32,
    parameter CHANNELS = 3,
    parameter FILTERS  = 28,
    parameter K        = 3,
    parameter PAD      = 1
)(
    input  wire clk,
    input  wire rst,
    input  wire start,
    output reg  done
);

    //--------------------------------------------------
    // Memories (NO file I/O here)
    //--------------------------------------------------
    reg [7:0] image_r [0:HEIGHT-1][0:WIDTH-1];
    reg [7:0] image_g [0:HEIGHT-1][0:WIDTH-1];
    reg [7:0] image_b [0:HEIGHT-1][0:WIDTH-1];

    reg signed [7:0] kernel [0:26][0:FILTERS-1];
    reg signed [7:0] bias   [0:FILTERS-1];

    reg signed [20:0] feature_map [0:FILTERS-1][0:HEIGHT-1][0:WIDTH-1];

    //--------------------------------------------------
    // Internal variables
    //--------------------------------------------------
    integer f,i,j,c,m,n;
    integer in_x,in_y,row_idx;

    reg signed [28:0] accum;
    reg signed [28:0] numerator;
    reg signed [23:0] kernel_mul;
    reg signed [23:0] bias_times_255;
    reg signed [20:0] out_int;
    reg signed [20:0] out_int_relu;

    reg [7:0] pix8;
    reg signed [15:0] kern16;
    reg signed [15:0] bias16;

    localparam IDLE=0, RUN=1, FIN=2;
    reg [1:0] state;

    //--------------------------------------------------
    // Sequential control
    //--------------------------------------------------
    always @(posedge clk or posedge rst) begin
        if(rst) begin
            state <= IDLE;
            done  <= 0;
        end
        else begin
            case(state)

            IDLE: begin
                done <= 0;
                if(start)
                    state <= RUN;
            end

            RUN: begin

                for(f=0; f<FILTERS; f=f+1) begin

                    bias16 = bias[f];
                    bias_times_255 = bias16 * 32'sd255;

                    for(i=0;i<HEIGHT;i=i+1) begin
                        for(j=0;j<WIDTH;j=j+1) begin

                            accum = bias_times_255;

                            for(m=0;m<K;m=m+1)
                                for(n=0;n<K;n=n+1) begin

                                    in_y = i + m - PAD;
                                    in_x = j + n - PAD;

                                    if(!(in_y<0 || in_y>=HEIGHT ||
                                         in_x<0 || in_x>=WIDTH)) begin

                                        for(c=0;c<CHANNELS;c=c+1) begin

                                            case(c)
                                                0: pix8 = image_r[in_y][in_x];
                                                1: pix8 = image_g[in_y][in_x];
                                                2: pix8 = image_b[in_y][in_x];
                                            endcase

                                            row_idx = m*K*CHANNELS + n*CHANNELS + c;
                                            kern16  = kernel[row_idx][f];

                                            // EXACT original multiply
                                            kernel_mul = kern16 * $signed({8'd0,pix8});
                                            accum = accum + kernel_mul;
                                        end
                                    end
                                end

                            numerator = accum;

                            // EXACT original rounding
                            if(numerator>=0)
                                out_int = (numerator + 32'sd127)/32'sd255;
                            else
                                out_int = -((-numerator + 32'sd127)/32'sd255);

                            if(out_int<0)
                                out_int_relu = 0;
                            else
                                out_int_relu = out_int;

                            feature_map[f][i][j] <= out_int_relu;
                        end
                    end
                end

                state <= FIN;
            end

            FIN: begin
                done <= 1;
                state <= IDLE;
            end

            endcase
        end
    end

endmodule
