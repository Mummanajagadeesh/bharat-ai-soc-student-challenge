module rom_07_conv2d_5_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:575][0:63];

    initial begin
        rom[0][0] = 8'd9;
        rom[0][1] = 8'd21;
        rom[0][2] = -8'd15;
        rom[0][3] = -8'd49;
        rom[0][4] = -8'd33;
        rom[0][5] = 8'd15;
        rom[0][6] = 8'd3;
        rom[0][7] = 8'd17;
        rom[0][8] = 8'd1;
        rom[0][9] = 8'd10;
        rom[0][10] = 8'd2;
        rom[0][11] = 8'd1;
        rom[0][12] = -8'd5;
        rom[0][13] = -8'd37;
        rom[0][14] = -8'd29;
        rom[0][15] = -8'd1;
        rom[0][16] = 8'd17;
        rom[0][17] = -8'd11;
        rom[0][18] = 8'd0;
        rom[0][19] = 8'd15;
        rom[0][20] = -8'd15;
        rom[0][21] = 8'd2;
        rom[0][22] = -8'd31;
        rom[0][23] = -8'd33;
        rom[0][24] = 8'd41;
        rom[0][25] = 8'd3;
        rom[0][26] = 8'd4;
        rom[0][27] = -8'd3;
        rom[0][28] = 8'd3;
        rom[0][29] = 8'd7;
        rom[0][30] = -8'd37;
        rom[0][31] = -8'd19;
        rom[0][32] = -8'd8;
        rom[0][33] = -8'd41;
        rom[0][34] = -8'd7;
        rom[0][35] = -8'd21;
        rom[0][36] = -8'd5;
        rom[0][37] = 8'd2;
        rom[0][38] = -8'd3;
        rom[0][39] = -8'd13;
        rom[0][40] = -8'd2;
        rom[0][41] = -8'd43;
        rom[0][42] = 8'd8;
        rom[0][43] = 8'd20;
        rom[0][44] = -8'd3;
        rom[0][45] = 8'd2;
        rom[0][46] = 8'd14;
        rom[0][47] = -8'd8;
        rom[0][48] = -8'd12;
        rom[0][49] = 8'd16;
        rom[0][50] = -8'd20;
        rom[0][51] = 8'd2;
        rom[0][52] = -8'd10;
        rom[0][53] = 8'd8;
        rom[0][54] = -8'd48;
        rom[0][55] = -8'd15;
        rom[0][56] = -8'd25;
        rom[0][57] = 8'd2;
        rom[0][58] = 8'd12;
        rom[0][59] = -8'd16;
        rom[0][60] = -8'd2;
        rom[0][61] = -8'd6;
        rom[0][62] = 8'd35;
        rom[0][63] = 8'd8;
        rom[1][0] = -8'd46;
        rom[1][1] = 8'd0;
        rom[1][2] = 8'd2;
        rom[1][3] = -8'd36;
        rom[1][4] = 8'd16;
        rom[1][5] = -8'd51;
        rom[1][6] = -8'd90;
        rom[1][7] = -8'd69;
        rom[1][8] = 8'd5;
        rom[1][9] = 8'd18;
        rom[1][10] = -8'd113;
        rom[1][11] = -8'd19;
        rom[1][12] = -8'd36;
        rom[1][13] = 8'd4;
        rom[1][14] = -8'd26;
        rom[1][15] = -8'd10;
        rom[1][16] = -8'd51;
        rom[1][17] = -8'd5;
        rom[1][18] = -8'd26;
        rom[1][19] = -8'd12;
        rom[1][20] = 8'd1;
        rom[1][21] = 8'd64;
        rom[1][22] = -8'd35;
        rom[1][23] = -8'd17;
        rom[1][24] = -8'd14;
        rom[1][25] = -8'd18;
        rom[1][26] = 8'd4;
        rom[1][27] = -8'd36;
        rom[1][28] = 8'd24;
        rom[1][29] = -8'd26;
        rom[1][30] = 8'd17;
        rom[1][31] = -8'd38;
        rom[1][32] = -8'd58;
        rom[1][33] = -8'd79;
        rom[1][34] = 8'd1;
        rom[1][35] = 8'd21;
        rom[1][36] = 8'd5;
        rom[1][37] = -8'd4;
        rom[1][38] = -8'd76;
        rom[1][39] = -8'd33;
        rom[1][40] = -8'd6;
        rom[1][41] = -8'd3;
        rom[1][42] = -8'd8;
        rom[1][43] = 8'd25;
        rom[1][44] = -8'd39;
        rom[1][45] = -8'd22;
        rom[1][46] = -8'd17;
        rom[1][47] = -8'd36;
        rom[1][48] = -8'd60;
        rom[1][49] = -8'd10;
        rom[1][50] = -8'd18;
        rom[1][51] = -8'd6;
        rom[1][52] = 8'd36;
        rom[1][53] = 8'd9;
        rom[1][54] = 8'd40;
        rom[1][55] = -8'd22;
        rom[1][56] = 8'd53;
        rom[1][57] = 8'd12;
        rom[1][58] = -8'd6;
        rom[1][59] = -8'd15;
        rom[1][60] = -8'd15;
        rom[1][61] = -8'd36;
        rom[1][62] = -8'd25;
        rom[1][63] = -8'd35;
        rom[2][0] = 8'd5;
        rom[2][1] = -8'd6;
        rom[2][2] = -8'd6;
        rom[2][3] = 8'd21;
        rom[2][4] = 8'd32;
        rom[2][5] = -8'd27;
        rom[2][6] = -8'd22;
        rom[2][7] = 8'd32;
        rom[2][8] = 8'd25;
        rom[2][9] = 8'd40;
        rom[2][10] = 8'd26;
        rom[2][11] = 8'd0;
        rom[2][12] = -8'd39;
        rom[2][13] = 8'd32;
        rom[2][14] = -8'd53;
        rom[2][15] = 8'd34;
        rom[2][16] = -8'd23;
        rom[2][17] = -8'd27;
        rom[2][18] = 8'd3;
        rom[2][19] = 8'd19;
        rom[2][20] = 8'd0;
        rom[2][21] = -8'd62;
        rom[2][22] = 8'd29;
        rom[2][23] = -8'd1;
        rom[2][24] = -8'd14;
        rom[2][25] = 8'd3;
        rom[2][26] = 8'd22;
        rom[2][27] = -8'd23;
        rom[2][28] = 8'd4;
        rom[2][29] = 8'd18;
        rom[2][30] = 8'd2;
        rom[2][31] = -8'd8;
        rom[2][32] = -8'd67;
        rom[2][33] = -8'd29;
        rom[2][34] = 8'd12;
        rom[2][35] = -8'd46;
        rom[2][36] = -8'd12;
        rom[2][37] = 8'd18;
        rom[2][38] = 8'd36;
        rom[2][39] = 8'd12;
        rom[2][40] = -8'd36;
        rom[2][41] = 8'd7;
        rom[2][42] = -8'd17;
        rom[2][43] = -8'd43;
        rom[2][44] = -8'd46;
        rom[2][45] = 8'd9;
        rom[2][46] = -8'd23;
        rom[2][47] = 8'd41;
        rom[2][48] = 8'd41;
        rom[2][49] = -8'd27;
        rom[2][50] = 8'd16;
        rom[2][51] = 8'd47;
        rom[2][52] = 8'd8;
        rom[2][53] = -8'd39;
        rom[2][54] = 8'd32;
        rom[2][55] = 8'd5;
        rom[2][56] = -8'd9;
        rom[2][57] = -8'd8;
        rom[2][58] = 8'd42;
        rom[2][59] = 8'd16;
        rom[2][60] = -8'd41;
        rom[2][61] = -8'd10;
        rom[2][62] = 8'd4;
        rom[2][63] = -8'd12;
        rom[3][0] = -8'd9;
        rom[3][1] = 8'd20;
        rom[3][2] = -8'd8;
        rom[3][3] = -8'd9;
        rom[3][4] = 8'd4;
        rom[3][5] = 8'd4;
        rom[3][6] = 8'd21;
        rom[3][7] = 8'd2;
        rom[3][8] = -8'd61;
        rom[3][9] = -8'd41;
        rom[3][10] = -8'd9;
        rom[3][11] = 8'd5;
        rom[3][12] = 8'd40;
        rom[3][13] = 8'd6;
        rom[3][14] = -8'd3;
        rom[3][15] = 8'd19;
        rom[3][16] = 8'd18;
        rom[3][17] = -8'd69;
        rom[3][18] = 8'd8;
        rom[3][19] = 8'd52;
        rom[3][20] = -8'd3;
        rom[3][21] = -8'd30;
        rom[3][22] = -8'd21;
        rom[3][23] = 8'd6;
        rom[3][24] = 8'd28;
        rom[3][25] = 8'd21;
        rom[3][26] = -8'd47;
        rom[3][27] = -8'd42;
        rom[3][28] = -8'd22;
        rom[3][29] = 8'd1;
        rom[3][30] = -8'd13;
        rom[3][31] = -8'd26;
        rom[3][32] = 8'd44;
        rom[3][33] = 8'd32;
        rom[3][34] = -8'd56;
        rom[3][35] = -8'd18;
        rom[3][36] = -8'd27;
        rom[3][37] = -8'd11;
        rom[3][38] = 8'd39;
        rom[3][39] = 8'd52;
        rom[3][40] = 8'd7;
        rom[3][41] = -8'd1;
        rom[3][42] = -8'd4;
        rom[3][43] = 8'd20;
        rom[3][44] = 8'd24;
        rom[3][45] = -8'd7;
        rom[3][46] = 8'd17;
        rom[3][47] = 8'd61;
        rom[3][48] = 8'd2;
        rom[3][49] = 8'd26;
        rom[3][50] = 8'd29;
        rom[3][51] = 8'd5;
        rom[3][52] = 8'd13;
        rom[3][53] = 8'd46;
        rom[3][54] = -8'd24;
        rom[3][55] = -8'd11;
        rom[3][56] = -8'd25;
        rom[3][57] = -8'd27;
        rom[3][58] = 8'd37;
        rom[3][59] = -8'd42;
        rom[3][60] = -8'd47;
        rom[3][61] = 8'd17;
        rom[3][62] = 8'd7;
        rom[3][63] = 8'd11;
        rom[4][0] = -8'd4;
        rom[4][1] = -8'd18;
        rom[4][2] = 8'd3;
        rom[4][3] = 8'd2;
        rom[4][4] = -8'd6;
        rom[4][5] = 8'd7;
        rom[4][6] = -8'd1;
        rom[4][7] = 8'd3;
        rom[4][8] = 8'd37;
        rom[4][9] = 8'd13;
        rom[4][10] = -8'd3;
        rom[4][11] = -8'd1;
        rom[4][12] = -8'd15;
        rom[4][13] = -8'd2;
        rom[4][14] = 8'd17;
        rom[4][15] = -8'd7;
        rom[4][16] = 8'd12;
        rom[4][17] = 8'd16;
        rom[4][18] = 8'd7;
        rom[4][19] = 8'd4;
        rom[4][20] = -8'd7;
        rom[4][21] = -8'd31;
        rom[4][22] = 8'd5;
        rom[4][23] = 8'd6;
        rom[4][24] = 8'd26;
        rom[4][25] = 8'd8;
        rom[4][26] = 8'd9;
        rom[4][27] = -8'd17;
        rom[4][28] = 8'd5;
        rom[4][29] = -8'd1;
        rom[4][30] = 8'd13;
        rom[4][31] = 8'd24;
        rom[4][32] = -8'd16;
        rom[4][33] = -8'd19;
        rom[4][34] = -8'd10;
        rom[4][35] = -8'd20;
        rom[4][36] = -8'd47;
        rom[4][37] = -8'd8;
        rom[4][38] = -8'd62;
        rom[4][39] = 8'd19;
        rom[4][40] = -8'd9;
        rom[4][41] = 8'd2;
        rom[4][42] = 8'd14;
        rom[4][43] = 8'd19;
        rom[4][44] = -8'd4;
        rom[4][45] = -8'd13;
        rom[4][46] = -8'd11;
        rom[4][47] = -8'd82;
        rom[4][48] = 8'd5;
        rom[4][49] = -8'd16;
        rom[4][50] = 8'd31;
        rom[4][51] = 8'd14;
        rom[4][52] = -8'd7;
        rom[4][53] = -8'd22;
        rom[4][54] = -8'd22;
        rom[4][55] = 8'd5;
        rom[4][56] = -8'd24;
        rom[4][57] = -8'd11;
        rom[4][58] = -8'd9;
        rom[4][59] = -8'd12;
        rom[4][60] = 8'd11;
        rom[4][61] = 8'd6;
        rom[4][62] = -8'd29;
        rom[4][63] = -8'd16;
        rom[5][0] = 8'd8;
        rom[5][1] = 8'd5;
        rom[5][2] = 8'd11;
        rom[5][3] = 8'd6;
        rom[5][4] = -8'd3;
        rom[5][5] = 8'd7;
        rom[5][6] = 8'd2;
        rom[5][7] = 8'd2;
        rom[5][8] = 8'd5;
        rom[5][9] = -8'd14;
        rom[5][10] = -8'd1;
        rom[5][11] = 8'd11;
        rom[5][12] = -8'd5;
        rom[5][13] = 8'd7;
        rom[5][14] = 8'd4;
        rom[5][15] = 8'd2;
        rom[5][16] = 8'd12;
        rom[5][17] = 8'd10;
        rom[5][18] = -8'd2;
        rom[5][19] = 8'd9;
        rom[5][20] = 8'd0;
        rom[5][21] = -8'd4;
        rom[5][22] = 8'd0;
        rom[5][23] = 8'd14;
        rom[5][24] = 8'd16;
        rom[5][25] = 8'd6;
        rom[5][26] = -8'd4;
        rom[5][27] = -8'd5;
        rom[5][28] = -8'd8;
        rom[5][29] = -8'd11;
        rom[5][30] = -8'd7;
        rom[5][31] = -8'd8;
        rom[5][32] = -8'd8;
        rom[5][33] = 8'd2;
        rom[5][34] = 8'd2;
        rom[5][35] = -8'd7;
        rom[5][36] = -8'd6;
        rom[5][37] = 8'd11;
        rom[5][38] = 8'd5;
        rom[5][39] = 8'd1;
        rom[5][40] = 8'd0;
        rom[5][41] = -8'd3;
        rom[5][42] = 8'd9;
        rom[5][43] = 8'd6;
        rom[5][44] = -8'd5;
        rom[5][45] = -8'd14;
        rom[5][46] = 8'd0;
        rom[5][47] = -8'd6;
        rom[5][48] = 8'd6;
        rom[5][49] = 8'd4;
        rom[5][50] = -8'd2;
        rom[5][51] = -8'd8;
        rom[5][52] = 8'd8;
        rom[5][53] = 8'd0;
        rom[5][54] = 8'd2;
        rom[5][55] = 8'd2;
        rom[5][56] = -8'd3;
        rom[5][57] = 8'd9;
        rom[5][58] = -8'd9;
        rom[5][59] = -8'd1;
        rom[5][60] = 8'd9;
        rom[5][61] = -8'd6;
        rom[5][62] = 8'd6;
        rom[5][63] = -8'd6;
        rom[6][0] = -8'd8;
        rom[6][1] = -8'd44;
        rom[6][2] = 8'd4;
        rom[6][3] = 8'd19;
        rom[6][4] = -8'd10;
        rom[6][5] = 8'd26;
        rom[6][6] = -8'd12;
        rom[6][7] = -8'd24;
        rom[6][8] = 8'd14;
        rom[6][9] = 8'd16;
        rom[6][10] = -8'd49;
        rom[6][11] = -8'd6;
        rom[6][12] = 8'd0;
        rom[6][13] = -8'd36;
        rom[6][14] = 8'd20;
        rom[6][15] = -8'd16;
        rom[6][16] = 8'd20;
        rom[6][17] = -8'd79;
        rom[6][18] = -8'd19;
        rom[6][19] = 8'd9;
        rom[6][20] = -8'd15;
        rom[6][21] = -8'd36;
        rom[6][22] = -8'd16;
        rom[6][23] = -8'd2;
        rom[6][24] = -8'd8;
        rom[6][25] = -8'd26;
        rom[6][26] = 8'd8;
        rom[6][27] = 8'd1;
        rom[6][28] = 8'd6;
        rom[6][29] = 8'd6;
        rom[6][30] = 8'd22;
        rom[6][31] = -8'd9;
        rom[6][32] = -8'd3;
        rom[6][33] = 8'd29;
        rom[6][34] = -8'd5;
        rom[6][35] = 8'd9;
        rom[6][36] = 8'd3;
        rom[6][37] = 8'd2;
        rom[6][38] = 8'd35;
        rom[6][39] = -8'd24;
        rom[6][40] = -8'd7;
        rom[6][41] = -8'd16;
        rom[6][42] = 8'd34;
        rom[6][43] = -8'd9;
        rom[6][44] = -8'd23;
        rom[6][45] = -8'd24;
        rom[6][46] = -8'd19;
        rom[6][47] = -8'd24;
        rom[6][48] = 8'd12;
        rom[6][49] = -8'd2;
        rom[6][50] = 8'd11;
        rom[6][51] = 8'd29;
        rom[6][52] = -8'd11;
        rom[6][53] = 8'd1;
        rom[6][54] = -8'd8;
        rom[6][55] = -8'd16;
        rom[6][56] = -8'd17;
        rom[6][57] = -8'd5;
        rom[6][58] = 8'd7;
        rom[6][59] = 8'd7;
        rom[6][60] = 8'd23;
        rom[6][61] = 8'd12;
        rom[6][62] = -8'd12;
        rom[6][63] = 8'd21;
        rom[7][0] = -8'd49;
        rom[7][1] = 8'd31;
        rom[7][2] = -8'd47;
        rom[7][3] = -8'd45;
        rom[7][4] = 8'd7;
        rom[7][5] = -8'd9;
        rom[7][6] = -8'd27;
        rom[7][7] = -8'd16;
        rom[7][8] = -8'd19;
        rom[7][9] = 8'd21;
        rom[7][10] = 8'd34;
        rom[7][11] = -8'd18;
        rom[7][12] = 8'd2;
        rom[7][13] = 8'd35;
        rom[7][14] = -8'd40;
        rom[7][15] = -8'd36;
        rom[7][16] = -8'd8;
        rom[7][17] = -8'd8;
        rom[7][18] = 8'd7;
        rom[7][19] = -8'd51;
        rom[7][20] = -8'd3;
        rom[7][21] = 8'd23;
        rom[7][22] = 8'd11;
        rom[7][23] = -8'd8;
        rom[7][24] = 8'd37;
        rom[7][25] = -8'd33;
        rom[7][26] = -8'd14;
        rom[7][27] = -8'd4;
        rom[7][28] = 8'd10;
        rom[7][29] = -8'd23;
        rom[7][30] = -8'd4;
        rom[7][31] = -8'd5;
        rom[7][32] = -8'd21;
        rom[7][33] = 8'd7;
        rom[7][34] = -8'd8;
        rom[7][35] = 8'd16;
        rom[7][36] = -8'd1;
        rom[7][37] = -8'd28;
        rom[7][38] = 8'd21;
        rom[7][39] = -8'd6;
        rom[7][40] = 8'd15;
        rom[7][41] = 8'd11;
        rom[7][42] = -8'd44;
        rom[7][43] = 8'd47;
        rom[7][44] = 8'd38;
        rom[7][45] = 8'd19;
        rom[7][46] = 8'd4;
        rom[7][47] = -8'd26;
        rom[7][48] = -8'd35;
        rom[7][49] = -8'd35;
        rom[7][50] = -8'd22;
        rom[7][51] = -8'd32;
        rom[7][52] = 8'd22;
        rom[7][53] = -8'd1;
        rom[7][54] = -8'd8;
        rom[7][55] = -8'd3;
        rom[7][56] = 8'd7;
        rom[7][57] = -8'd19;
        rom[7][58] = -8'd81;
        rom[7][59] = 8'd12;
        rom[7][60] = -8'd16;
        rom[7][61] = -8'd79;
        rom[7][62] = 8'd0;
        rom[7][63] = 8'd41;
        rom[8][0] = -8'd13;
        rom[8][1] = 8'd27;
        rom[8][2] = -8'd11;
        rom[8][3] = 8'd16;
        rom[8][4] = -8'd13;
        rom[8][5] = -8'd6;
        rom[8][6] = 8'd9;
        rom[8][7] = 8'd33;
        rom[8][8] = 8'd0;
        rom[8][9] = 8'd29;
        rom[8][10] = -8'd4;
        rom[8][11] = -8'd22;
        rom[8][12] = 8'd10;
        rom[8][13] = 8'd18;
        rom[8][14] = 8'd6;
        rom[8][15] = 8'd47;
        rom[8][16] = 8'd6;
        rom[8][17] = 8'd6;
        rom[8][18] = -8'd18;
        rom[8][19] = 8'd22;
        rom[8][20] = -8'd1;
        rom[8][21] = 8'd13;
        rom[8][22] = -8'd18;
        rom[8][23] = -8'd7;
        rom[8][24] = 8'd16;
        rom[8][25] = 8'd2;
        rom[8][26] = -8'd19;
        rom[8][27] = -8'd42;
        rom[8][28] = 8'd5;
        rom[8][29] = -8'd30;
        rom[8][30] = 8'd14;
        rom[8][31] = 8'd20;
        rom[8][32] = 8'd0;
        rom[8][33] = -8'd38;
        rom[8][34] = -8'd3;
        rom[8][35] = -8'd23;
        rom[8][36] = -8'd19;
        rom[8][37] = 8'd11;
        rom[8][38] = -8'd24;
        rom[8][39] = -8'd18;
        rom[8][40] = -8'd29;
        rom[8][41] = 8'd6;
        rom[8][42] = 8'd2;
        rom[8][43] = 8'd5;
        rom[8][44] = -8'd11;
        rom[8][45] = -8'd3;
        rom[8][46] = 8'd34;
        rom[8][47] = 8'd19;
        rom[8][48] = -8'd22;
        rom[8][49] = -8'd48;
        rom[8][50] = 8'd11;
        rom[8][51] = 8'd6;
        rom[8][52] = 8'd5;
        rom[8][53] = 8'd11;
        rom[8][54] = 8'd13;
        rom[8][55] = 8'd3;
        rom[8][56] = -8'd38;
        rom[8][57] = -8'd7;
        rom[8][58] = 8'd27;
        rom[8][59] = -8'd1;
        rom[8][60] = 8'd4;
        rom[8][61] = -8'd64;
        rom[8][62] = -8'd25;
        rom[8][63] = -8'd26;
        rom[9][0] = 8'd6;
        rom[9][1] = 8'd28;
        rom[9][2] = 8'd2;
        rom[9][3] = -8'd50;
        rom[9][4] = 8'd15;
        rom[9][5] = 8'd3;
        rom[9][6] = 8'd19;
        rom[9][7] = 8'd1;
        rom[9][8] = -8'd20;
        rom[9][9] = 8'd14;
        rom[9][10] = 8'd5;
        rom[9][11] = -8'd30;
        rom[9][12] = -8'd17;
        rom[9][13] = 8'd15;
        rom[9][14] = 8'd11;
        rom[9][15] = -8'd26;
        rom[9][16] = 8'd15;
        rom[9][17] = 8'd6;
        rom[9][18] = 8'd20;
        rom[9][19] = -8'd70;
        rom[9][20] = -8'd13;
        rom[9][21] = 8'd16;
        rom[9][22] = -8'd42;
        rom[9][23] = 8'd22;
        rom[9][24] = 8'd30;
        rom[9][25] = -8'd13;
        rom[9][26] = -8'd7;
        rom[9][27] = -8'd27;
        rom[9][28] = -8'd33;
        rom[9][29] = 8'd24;
        rom[9][30] = 8'd3;
        rom[9][31] = 8'd12;
        rom[9][32] = 8'd22;
        rom[9][33] = -8'd1;
        rom[9][34] = -8'd2;
        rom[9][35] = -8'd20;
        rom[9][36] = 8'd26;
        rom[9][37] = 8'd55;
        rom[9][38] = 8'd31;
        rom[9][39] = -8'd29;
        rom[9][40] = -8'd11;
        rom[9][41] = 8'd10;
        rom[9][42] = -8'd48;
        rom[9][43] = -8'd31;
        rom[9][44] = -8'd18;
        rom[9][45] = -8'd22;
        rom[9][46] = -8'd17;
        rom[9][47] = -8'd23;
        rom[9][48] = -8'd17;
        rom[9][49] = 8'd12;
        rom[9][50] = -8'd47;
        rom[9][51] = 8'd14;
        rom[9][52] = 8'd26;
        rom[9][53] = -8'd3;
        rom[9][54] = -8'd23;
        rom[9][55] = 8'd20;
        rom[9][56] = 8'd5;
        rom[9][57] = -8'd52;
        rom[9][58] = -8'd41;
        rom[9][59] = -8'd9;
        rom[9][60] = 8'd27;
        rom[9][61] = -8'd7;
        rom[9][62] = 8'd18;
        rom[9][63] = -8'd7;
        rom[10][0] = 8'd0;
        rom[10][1] = 8'd32;
        rom[10][2] = 8'd18;
        rom[10][3] = 8'd4;
        rom[10][4] = -8'd19;
        rom[10][5] = 8'd11;
        rom[10][6] = 8'd49;
        rom[10][7] = -8'd10;
        rom[10][8] = 8'd25;
        rom[10][9] = 8'd19;
        rom[10][10] = 8'd3;
        rom[10][11] = 8'd26;
        rom[10][12] = -8'd24;
        rom[10][13] = -8'd36;
        rom[10][14] = -8'd14;
        rom[10][15] = -8'd11;
        rom[10][16] = -8'd8;
        rom[10][17] = -8'd37;
        rom[10][18] = 8'd0;
        rom[10][19] = -8'd23;
        rom[10][20] = -8'd2;
        rom[10][21] = -8'd11;
        rom[10][22] = -8'd25;
        rom[10][23] = -8'd30;
        rom[10][24] = -8'd9;
        rom[10][25] = -8'd128;
        rom[10][26] = 8'd21;
        rom[10][27] = 8'd8;
        rom[10][28] = -8'd41;
        rom[10][29] = 8'd13;
        rom[10][30] = -8'd3;
        rom[10][31] = 8'd38;
        rom[10][32] = 8'd26;
        rom[10][33] = 8'd15;
        rom[10][34] = -8'd75;
        rom[10][35] = -8'd18;
        rom[10][36] = 8'd46;
        rom[10][37] = 8'd31;
        rom[10][38] = 8'd50;
        rom[10][39] = 8'd21;
        rom[10][40] = 8'd10;
        rom[10][41] = -8'd15;
        rom[10][42] = -8'd18;
        rom[10][43] = -8'd20;
        rom[10][44] = -8'd26;
        rom[10][45] = -8'd12;
        rom[10][46] = 8'd13;
        rom[10][47] = 8'd10;
        rom[10][48] = 8'd18;
        rom[10][49] = 8'd4;
        rom[10][50] = -8'd19;
        rom[10][51] = 8'd3;
        rom[10][52] = -8'd1;
        rom[10][53] = -8'd93;
        rom[10][54] = -8'd20;
        rom[10][55] = -8'd15;
        rom[10][56] = 8'd29;
        rom[10][57] = 8'd40;
        rom[10][58] = 8'd16;
        rom[10][59] = 8'd11;
        rom[10][60] = -8'd1;
        rom[10][61] = -8'd29;
        rom[10][62] = 8'd1;
        rom[10][63] = -8'd3;
        rom[11][0] = 8'd35;
        rom[11][1] = 8'd33;
        rom[11][2] = 8'd15;
        rom[11][3] = -8'd32;
        rom[11][4] = 8'd7;
        rom[11][5] = 8'd20;
        rom[11][6] = -8'd7;
        rom[11][7] = 8'd38;
        rom[11][8] = 8'd29;
        rom[11][9] = -8'd43;
        rom[11][10] = 8'd4;
        rom[11][11] = -8'd17;
        rom[11][12] = -8'd6;
        rom[11][13] = -8'd22;
        rom[11][14] = 8'd29;
        rom[11][15] = 8'd28;
        rom[11][16] = -8'd20;
        rom[11][17] = 8'd56;
        rom[11][18] = -8'd28;
        rom[11][19] = -8'd3;
        rom[11][20] = -8'd11;
        rom[11][21] = -8'd25;
        rom[11][22] = 8'd57;
        rom[11][23] = 8'd0;
        rom[11][24] = 8'd0;
        rom[11][25] = 8'd18;
        rom[11][26] = 8'd6;
        rom[11][27] = 8'd21;
        rom[11][28] = -8'd31;
        rom[11][29] = 8'd4;
        rom[11][30] = -8'd23;
        rom[11][31] = 8'd57;
        rom[11][32] = -8'd34;
        rom[11][33] = 8'd12;
        rom[11][34] = -8'd1;
        rom[11][35] = -8'd4;
        rom[11][36] = 8'd18;
        rom[11][37] = 8'd5;
        rom[11][38] = 8'd19;
        rom[11][39] = -8'd41;
        rom[11][40] = 8'd24;
        rom[11][41] = 8'd23;
        rom[11][42] = -8'd24;
        rom[11][43] = 8'd19;
        rom[11][44] = 8'd29;
        rom[11][45] = 8'd28;
        rom[11][46] = -8'd10;
        rom[11][47] = 8'd1;
        rom[11][48] = 8'd12;
        rom[11][49] = -8'd1;
        rom[11][50] = -8'd14;
        rom[11][51] = -8'd38;
        rom[11][52] = 8'd0;
        rom[11][53] = 8'd2;
        rom[11][54] = 8'd47;
        rom[11][55] = 8'd54;
        rom[11][56] = 8'd10;
        rom[11][57] = -8'd22;
        rom[11][58] = -8'd24;
        rom[11][59] = -8'd16;
        rom[11][60] = 8'd23;
        rom[11][61] = 8'd29;
        rom[11][62] = -8'd25;
        rom[11][63] = 8'd43;
        rom[12][0] = 8'd5;
        rom[12][1] = 8'd4;
        rom[12][2] = 8'd48;
        rom[12][3] = -8'd42;
        rom[12][4] = -8'd35;
        rom[12][5] = -8'd7;
        rom[12][6] = 8'd5;
        rom[12][7] = 8'd44;
        rom[12][8] = 8'd11;
        rom[12][9] = 8'd19;
        rom[12][10] = 8'd10;
        rom[12][11] = 8'd39;
        rom[12][12] = -8'd37;
        rom[12][13] = 8'd36;
        rom[12][14] = 8'd21;
        rom[12][15] = -8'd62;
        rom[12][16] = -8'd45;
        rom[12][17] = 8'd4;
        rom[12][18] = -8'd24;
        rom[12][19] = -8'd3;
        rom[12][20] = 8'd8;
        rom[12][21] = 8'd6;
        rom[12][22] = 8'd10;
        rom[12][23] = -8'd32;
        rom[12][24] = -8'd16;
        rom[12][25] = 8'd29;
        rom[12][26] = 8'd13;
        rom[12][27] = 8'd7;
        rom[12][28] = 8'd30;
        rom[12][29] = 8'd17;
        rom[12][30] = 8'd36;
        rom[12][31] = -8'd2;
        rom[12][32] = -8'd15;
        rom[12][33] = -8'd37;
        rom[12][34] = 8'd17;
        rom[12][35] = -8'd30;
        rom[12][36] = 8'd60;
        rom[12][37] = 8'd6;
        rom[12][38] = 8'd20;
        rom[12][39] = 8'd32;
        rom[12][40] = -8'd29;
        rom[12][41] = -8'd48;
        rom[12][42] = -8'd18;
        rom[12][43] = -8'd10;
        rom[12][44] = 8'd0;
        rom[12][45] = 8'd41;
        rom[12][46] = -8'd24;
        rom[12][47] = -8'd29;
        rom[12][48] = 8'd31;
        rom[12][49] = 8'd17;
        rom[12][50] = 8'd23;
        rom[12][51] = 8'd0;
        rom[12][52] = -8'd2;
        rom[12][53] = -8'd24;
        rom[12][54] = 8'd40;
        rom[12][55] = -8'd3;
        rom[12][56] = 8'd18;
        rom[12][57] = 8'd2;
        rom[12][58] = 8'd2;
        rom[12][59] = -8'd17;
        rom[12][60] = -8'd8;
        rom[12][61] = 8'd6;
        rom[12][62] = 8'd17;
        rom[12][63] = 8'd34;
        rom[13][0] = -8'd8;
        rom[13][1] = -8'd30;
        rom[13][2] = -8'd20;
        rom[13][3] = -8'd37;
        rom[13][4] = 8'd15;
        rom[13][5] = 8'd17;
        rom[13][6] = 8'd22;
        rom[13][7] = -8'd4;
        rom[13][8] = 8'd35;
        rom[13][9] = -8'd11;
        rom[13][10] = -8'd22;
        rom[13][11] = -8'd3;
        rom[13][12] = -8'd8;
        rom[13][13] = -8'd2;
        rom[13][14] = -8'd23;
        rom[13][15] = -8'd10;
        rom[13][16] = -8'd18;
        rom[13][17] = -8'd33;
        rom[13][18] = -8'd23;
        rom[13][19] = -8'd22;
        rom[13][20] = -8'd3;
        rom[13][21] = -8'd6;
        rom[13][22] = 8'd2;
        rom[13][23] = 8'd2;
        rom[13][24] = -8'd2;
        rom[13][25] = -8'd41;
        rom[13][26] = -8'd9;
        rom[13][27] = 8'd12;
        rom[13][28] = -8'd1;
        rom[13][29] = -8'd24;
        rom[13][30] = -8'd67;
        rom[13][31] = 8'd2;
        rom[13][32] = 8'd20;
        rom[13][33] = -8'd39;
        rom[13][34] = -8'd54;
        rom[13][35] = -8'd1;
        rom[13][36] = -8'd10;
        rom[13][37] = -8'd12;
        rom[13][38] = -8'd12;
        rom[13][39] = 8'd30;
        rom[13][40] = -8'd4;
        rom[13][41] = -8'd3;
        rom[13][42] = 8'd4;
        rom[13][43] = -8'd14;
        rom[13][44] = -8'd24;
        rom[13][45] = 8'd41;
        rom[13][46] = 8'd32;
        rom[13][47] = -8'd11;
        rom[13][48] = -8'd5;
        rom[13][49] = -8'd53;
        rom[13][50] = -8'd2;
        rom[13][51] = 8'd12;
        rom[13][52] = 8'd22;
        rom[13][53] = -8'd50;
        rom[13][54] = -8'd33;
        rom[13][55] = 8'd1;
        rom[13][56] = -8'd4;
        rom[13][57] = 8'd13;
        rom[13][58] = -8'd4;
        rom[13][59] = -8'd52;
        rom[13][60] = -8'd29;
        rom[13][61] = -8'd31;
        rom[13][62] = -8'd36;
        rom[13][63] = 8'd41;
        rom[14][0] = 8'd16;
        rom[14][1] = 8'd11;
        rom[14][2] = 8'd16;
        rom[14][3] = -8'd5;
        rom[14][4] = -8'd13;
        rom[14][5] = 8'd6;
        rom[14][6] = -8'd25;
        rom[14][7] = -8'd8;
        rom[14][8] = -8'd11;
        rom[14][9] = -8'd51;
        rom[14][10] = 8'd28;
        rom[14][11] = 8'd40;
        rom[14][12] = -8'd5;
        rom[14][13] = -8'd19;
        rom[14][14] = 8'd6;
        rom[14][15] = -8'd8;
        rom[14][16] = 8'd2;
        rom[14][17] = 8'd32;
        rom[14][18] = 8'd17;
        rom[14][19] = 8'd8;
        rom[14][20] = -8'd4;
        rom[14][21] = 8'd16;
        rom[14][22] = -8'd2;
        rom[14][23] = 8'd0;
        rom[14][24] = -8'd27;
        rom[14][25] = 8'd3;
        rom[14][26] = -8'd12;
        rom[14][27] = 8'd13;
        rom[14][28] = -8'd27;
        rom[14][29] = -8'd81;
        rom[14][30] = 8'd17;
        rom[14][31] = 8'd32;
        rom[14][32] = 8'd22;
        rom[14][33] = 8'd8;
        rom[14][34] = -8'd16;
        rom[14][35] = -8'd16;
        rom[14][36] = -8'd23;
        rom[14][37] = -8'd32;
        rom[14][38] = -8'd23;
        rom[14][39] = -8'd1;
        rom[14][40] = 8'd12;
        rom[14][41] = 8'd18;
        rom[14][42] = -8'd3;
        rom[14][43] = -8'd6;
        rom[14][44] = 8'd4;
        rom[14][45] = 8'd24;
        rom[14][46] = -8'd2;
        rom[14][47] = -8'd33;
        rom[14][48] = 8'd4;
        rom[14][49] = -8'd40;
        rom[14][50] = 8'd24;
        rom[14][51] = -8'd48;
        rom[14][52] = 8'd14;
        rom[14][53] = 8'd22;
        rom[14][54] = -8'd6;
        rom[14][55] = -8'd46;
        rom[14][56] = 8'd9;
        rom[14][57] = 8'd0;
        rom[14][58] = -8'd3;
        rom[14][59] = -8'd6;
        rom[14][60] = -8'd12;
        rom[14][61] = 8'd44;
        rom[14][62] = 8'd6;
        rom[14][63] = 8'd11;
        rom[15][0] = 8'd14;
        rom[15][1] = -8'd57;
        rom[15][2] = -8'd34;
        rom[15][3] = -8'd45;
        rom[15][4] = -8'd61;
        rom[15][5] = 8'd17;
        rom[15][6] = -8'd37;
        rom[15][7] = 8'd4;
        rom[15][8] = -8'd98;
        rom[15][9] = 8'd1;
        rom[15][10] = -8'd44;
        rom[15][11] = -8'd12;
        rom[15][12] = 8'd29;
        rom[15][13] = 8'd16;
        rom[15][14] = 8'd11;
        rom[15][15] = -8'd8;
        rom[15][16] = -8'd14;
        rom[15][17] = 8'd44;
        rom[15][18] = 8'd18;
        rom[15][19] = 8'd1;
        rom[15][20] = -8'd6;
        rom[15][21] = 8'd34;
        rom[15][22] = -8'd59;
        rom[15][23] = 8'd7;
        rom[15][24] = 8'd32;
        rom[15][25] = 8'd8;
        rom[15][26] = -8'd15;
        rom[15][27] = -8'd11;
        rom[15][28] = -8'd23;
        rom[15][29] = -8'd1;
        rom[15][30] = -8'd1;
        rom[15][31] = -8'd5;
        rom[15][32] = 8'd47;
        rom[15][33] = 8'd42;
        rom[15][34] = 8'd27;
        rom[15][35] = -8'd4;
        rom[15][36] = 8'd28;
        rom[15][37] = 8'd3;
        rom[15][38] = -8'd5;
        rom[15][39] = 8'd13;
        rom[15][40] = -8'd44;
        rom[15][41] = 8'd25;
        rom[15][42] = -8'd2;
        rom[15][43] = -8'd61;
        rom[15][44] = -8'd26;
        rom[15][45] = -8'd22;
        rom[15][46] = 8'd0;
        rom[15][47] = -8'd13;
        rom[15][48] = 8'd2;
        rom[15][49] = -8'd32;
        rom[15][50] = 8'd54;
        rom[15][51] = -8'd24;
        rom[15][52] = 8'd21;
        rom[15][53] = 8'd8;
        rom[15][54] = 8'd28;
        rom[15][55] = -8'd50;
        rom[15][56] = -8'd10;
        rom[15][57] = 8'd27;
        rom[15][58] = 8'd17;
        rom[15][59] = -8'd6;
        rom[15][60] = -8'd19;
        rom[15][61] = 8'd26;
        rom[15][62] = -8'd12;
        rom[15][63] = -8'd6;
        rom[16][0] = -8'd3;
        rom[16][1] = 8'd8;
        rom[16][2] = -8'd1;
        rom[16][3] = -8'd7;
        rom[16][4] = -8'd6;
        rom[16][5] = -8'd8;
        rom[16][6] = -8'd8;
        rom[16][7] = 8'd2;
        rom[16][8] = -8'd6;
        rom[16][9] = 8'd1;
        rom[16][10] = -8'd2;
        rom[16][11] = -8'd8;
        rom[16][12] = 8'd4;
        rom[16][13] = -8'd2;
        rom[16][14] = 8'd7;
        rom[16][15] = 8'd7;
        rom[16][16] = -8'd8;
        rom[16][17] = -8'd1;
        rom[16][18] = 8'd2;
        rom[16][19] = 8'd5;
        rom[16][20] = 8'd7;
        rom[16][21] = 8'd8;
        rom[16][22] = -8'd5;
        rom[16][23] = 8'd7;
        rom[16][24] = 8'd3;
        rom[16][25] = -8'd1;
        rom[16][26] = -8'd8;
        rom[16][27] = 8'd1;
        rom[16][28] = 8'd0;
        rom[16][29] = -8'd4;
        rom[16][30] = 8'd7;
        rom[16][31] = 8'd2;
        rom[16][32] = 8'd9;
        rom[16][33] = 8'd10;
        rom[16][34] = -8'd2;
        rom[16][35] = 8'd2;
        rom[16][36] = 8'd8;
        rom[16][37] = -8'd6;
        rom[16][38] = 8'd5;
        rom[16][39] = -8'd1;
        rom[16][40] = 8'd8;
        rom[16][41] = -8'd6;
        rom[16][42] = -8'd8;
        rom[16][43] = -8'd6;
        rom[16][44] = 8'd5;
        rom[16][45] = 8'd9;
        rom[16][46] = -8'd4;
        rom[16][47] = -8'd3;
        rom[16][48] = -8'd8;
        rom[16][49] = -8'd8;
        rom[16][50] = 8'd4;
        rom[16][51] = 8'd6;
        rom[16][52] = 8'd5;
        rom[16][53] = 8'd2;
        rom[16][54] = -8'd2;
        rom[16][55] = 8'd6;
        rom[16][56] = 8'd2;
        rom[16][57] = 8'd3;
        rom[16][58] = 8'd3;
        rom[16][59] = -8'd1;
        rom[16][60] = 8'd5;
        rom[16][61] = -8'd7;
        rom[16][62] = 8'd1;
        rom[16][63] = 8'd8;
        rom[17][0] = 8'd28;
        rom[17][1] = 8'd4;
        rom[17][2] = -8'd4;
        rom[17][3] = 8'd60;
        rom[17][4] = 8'd21;
        rom[17][5] = 8'd48;
        rom[17][6] = 8'd41;
        rom[17][7] = 8'd44;
        rom[17][8] = 8'd17;
        rom[17][9] = -8'd22;
        rom[17][10] = 8'd7;
        rom[17][11] = 8'd14;
        rom[17][12] = -8'd33;
        rom[17][13] = 8'd30;
        rom[17][14] = 8'd10;
        rom[17][15] = 8'd31;
        rom[17][16] = 8'd9;
        rom[17][17] = -8'd6;
        rom[17][18] = 8'd28;
        rom[17][19] = 8'd9;
        rom[17][20] = -8'd9;
        rom[17][21] = -8'd25;
        rom[17][22] = 8'd15;
        rom[17][23] = -8'd20;
        rom[17][24] = 8'd53;
        rom[17][25] = -8'd3;
        rom[17][26] = -8'd25;
        rom[17][27] = -8'd10;
        rom[17][28] = -8'd40;
        rom[17][29] = 8'd14;
        rom[17][30] = 8'd31;
        rom[17][31] = 8'd28;
        rom[17][32] = -8'd22;
        rom[17][33] = -8'd12;
        rom[17][34] = 8'd19;
        rom[17][35] = -8'd30;
        rom[17][36] = -8'd17;
        rom[17][37] = 8'd15;
        rom[17][38] = 8'd36;
        rom[17][39] = -8'd19;
        rom[17][40] = 8'd22;
        rom[17][41] = 8'd16;
        rom[17][42] = -8'd23;
        rom[17][43] = 8'd18;
        rom[17][44] = -8'd37;
        rom[17][45] = -8'd4;
        rom[17][46] = -8'd21;
        rom[17][47] = 8'd12;
        rom[17][48] = -8'd26;
        rom[17][49] = 8'd15;
        rom[17][50] = 8'd26;
        rom[17][51] = -8'd71;
        rom[17][52] = -8'd20;
        rom[17][53] = -8'd6;
        rom[17][54] = 8'd26;
        rom[17][55] = -8'd10;
        rom[17][56] = -8'd11;
        rom[17][57] = -8'd33;
        rom[17][58] = -8'd14;
        rom[17][59] = -8'd21;
        rom[17][60] = 8'd0;
        rom[17][61] = -8'd74;
        rom[17][62] = -8'd37;
        rom[17][63] = 8'd5;
        rom[18][0] = -8'd57;
        rom[18][1] = 8'd30;
        rom[18][2] = -8'd9;
        rom[18][3] = 8'd1;
        rom[18][4] = -8'd22;
        rom[18][5] = -8'd28;
        rom[18][6] = 8'd2;
        rom[18][7] = 8'd25;
        rom[18][8] = 8'd9;
        rom[18][9] = 8'd14;
        rom[18][10] = 8'd39;
        rom[18][11] = -8'd5;
        rom[18][12] = -8'd32;
        rom[18][13] = 8'd8;
        rom[18][14] = -8'd22;
        rom[18][15] = 8'd12;
        rom[18][16] = -8'd4;
        rom[18][17] = 8'd43;
        rom[18][18] = -8'd37;
        rom[18][19] = -8'd29;
        rom[18][20] = -8'd8;
        rom[18][21] = -8'd3;
        rom[18][22] = 8'd19;
        rom[18][23] = -8'd21;
        rom[18][24] = 8'd16;
        rom[18][25] = 8'd4;
        rom[18][26] = -8'd83;
        rom[18][27] = 8'd30;
        rom[18][28] = 8'd20;
        rom[18][29] = -8'd17;
        rom[18][30] = -8'd9;
        rom[18][31] = 8'd36;
        rom[18][32] = -8'd23;
        rom[18][33] = 8'd4;
        rom[18][34] = -8'd12;
        rom[18][35] = -8'd20;
        rom[18][36] = -8'd19;
        rom[18][37] = 8'd1;
        rom[18][38] = -8'd5;
        rom[18][39] = 8'd33;
        rom[18][40] = -8'd5;
        rom[18][41] = 8'd12;
        rom[18][42] = -8'd60;
        rom[18][43] = -8'd42;
        rom[18][44] = 8'd18;
        rom[18][45] = 8'd28;
        rom[18][46] = 8'd4;
        rom[18][47] = 8'd5;
        rom[18][48] = -8'd28;
        rom[18][49] = -8'd12;
        rom[18][50] = -8'd16;
        rom[18][51] = 8'd4;
        rom[18][52] = -8'd31;
        rom[18][53] = -8'd32;
        rom[18][54] = -8'd32;
        rom[18][55] = 8'd2;
        rom[18][56] = -8'd1;
        rom[18][57] = -8'd59;
        rom[18][58] = 8'd4;
        rom[18][59] = 8'd9;
        rom[18][60] = -8'd9;
        rom[18][61] = -8'd17;
        rom[18][62] = -8'd44;
        rom[18][63] = 8'd14;
        rom[19][0] = -8'd52;
        rom[19][1] = 8'd13;
        rom[19][2] = -8'd57;
        rom[19][3] = -8'd9;
        rom[19][4] = -8'd65;
        rom[19][5] = 8'd20;
        rom[19][6] = -8'd31;
        rom[19][7] = -8'd7;
        rom[19][8] = -8'd28;
        rom[19][9] = 8'd32;
        rom[19][10] = 8'd15;
        rom[19][11] = -8'd8;
        rom[19][12] = -8'd20;
        rom[19][13] = -8'd33;
        rom[19][14] = 8'd4;
        rom[19][15] = 8'd25;
        rom[19][16] = -8'd28;
        rom[19][17] = -8'd3;
        rom[19][18] = 8'd6;
        rom[19][19] = -8'd25;
        rom[19][20] = 8'd0;
        rom[19][21] = 8'd6;
        rom[19][22] = 8'd2;
        rom[19][23] = -8'd60;
        rom[19][24] = 8'd9;
        rom[19][25] = -8'd8;
        rom[19][26] = -8'd11;
        rom[19][27] = -8'd66;
        rom[19][28] = 8'd38;
        rom[19][29] = 8'd14;
        rom[19][30] = 8'd22;
        rom[19][31] = 8'd16;
        rom[19][32] = -8'd14;
        rom[19][33] = -8'd28;
        rom[19][34] = 8'd18;
        rom[19][35] = 8'd7;
        rom[19][36] = -8'd12;
        rom[19][37] = 8'd3;
        rom[19][38] = -8'd35;
        rom[19][39] = -8'd32;
        rom[19][40] = -8'd34;
        rom[19][41] = 8'd7;
        rom[19][42] = -8'd58;
        rom[19][43] = -8'd51;
        rom[19][44] = 8'd4;
        rom[19][45] = -8'd46;
        rom[19][46] = 8'd2;
        rom[19][47] = 8'd32;
        rom[19][48] = 8'd24;
        rom[19][49] = -8'd19;
        rom[19][50] = -8'd8;
        rom[19][51] = -8'd16;
        rom[19][52] = 8'd24;
        rom[19][53] = 8'd2;
        rom[19][54] = 8'd26;
        rom[19][55] = 8'd3;
        rom[19][56] = 8'd25;
        rom[19][57] = 8'd0;
        rom[19][58] = -8'd15;
        rom[19][59] = 8'd36;
        rom[19][60] = -8'd9;
        rom[19][61] = 8'd0;
        rom[19][62] = 8'd21;
        rom[19][63] = 8'd49;
        rom[20][0] = 8'd27;
        rom[20][1] = -8'd33;
        rom[20][2] = -8'd6;
        rom[20][3] = -8'd5;
        rom[20][4] = 8'd17;
        rom[20][5] = -8'd1;
        rom[20][6] = -8'd1;
        rom[20][7] = -8'd24;
        rom[20][8] = -8'd6;
        rom[20][9] = 8'd21;
        rom[20][10] = -8'd15;
        rom[20][11] = -8'd15;
        rom[20][12] = -8'd16;
        rom[20][13] = -8'd39;
        rom[20][14] = 8'd13;
        rom[20][15] = 8'd14;
        rom[20][16] = -8'd69;
        rom[20][17] = 8'd0;
        rom[20][18] = -8'd54;
        rom[20][19] = 8'd0;
        rom[20][20] = -8'd8;
        rom[20][21] = 8'd4;
        rom[20][22] = -8'd18;
        rom[20][23] = -8'd18;
        rom[20][24] = 8'd27;
        rom[20][25] = -8'd26;
        rom[20][26] = -8'd7;
        rom[20][27] = -8'd4;
        rom[20][28] = 8'd23;
        rom[20][29] = -8'd5;
        rom[20][30] = 8'd10;
        rom[20][31] = 8'd32;
        rom[20][32] = -8'd19;
        rom[20][33] = -8'd29;
        rom[20][34] = -8'd67;
        rom[20][35] = -8'd6;
        rom[20][36] = -8'd12;
        rom[20][37] = 8'd17;
        rom[20][38] = -8'd29;
        rom[20][39] = -8'd15;
        rom[20][40] = -8'd35;
        rom[20][41] = -8'd56;
        rom[20][42] = -8'd25;
        rom[20][43] = 8'd2;
        rom[20][44] = -8'd22;
        rom[20][45] = 8'd0;
        rom[20][46] = -8'd30;
        rom[20][47] = 8'd14;
        rom[20][48] = 8'd7;
        rom[20][49] = -8'd14;
        rom[20][50] = 8'd14;
        rom[20][51] = -8'd5;
        rom[20][52] = 8'd34;
        rom[20][53] = 8'd5;
        rom[20][54] = -8'd23;
        rom[20][55] = 8'd5;
        rom[20][56] = -8'd27;
        rom[20][57] = -8'd27;
        rom[20][58] = 8'd28;
        rom[20][59] = 8'd8;
        rom[20][60] = 8'd22;
        rom[20][61] = 8'd5;
        rom[20][62] = 8'd8;
        rom[20][63] = -8'd7;
        rom[21][0] = 8'd5;
        rom[21][1] = 8'd1;
        rom[21][2] = 8'd7;
        rom[21][3] = 8'd9;
        rom[21][4] = 8'd2;
        rom[21][5] = -8'd3;
        rom[21][6] = -8'd4;
        rom[21][7] = -8'd3;
        rom[21][8] = -8'd7;
        rom[21][9] = -8'd4;
        rom[21][10] = 8'd2;
        rom[21][11] = -8'd9;
        rom[21][12] = 8'd0;
        rom[21][13] = 8'd9;
        rom[21][14] = 8'd7;
        rom[21][15] = -8'd8;
        rom[21][16] = 8'd5;
        rom[21][17] = 8'd8;
        rom[21][18] = -8'd6;
        rom[21][19] = 8'd1;
        rom[21][20] = 8'd4;
        rom[21][21] = -8'd5;
        rom[21][22] = -8'd10;
        rom[21][23] = -8'd7;
        rom[21][24] = -8'd8;
        rom[21][25] = -8'd6;
        rom[21][26] = 8'd5;
        rom[21][27] = 8'd4;
        rom[21][28] = 8'd1;
        rom[21][29] = 8'd5;
        rom[21][30] = 8'd6;
        rom[21][31] = -8'd7;
        rom[21][32] = -8'd4;
        rom[21][33] = 8'd7;
        rom[21][34] = 8'd7;
        rom[21][35] = 8'd0;
        rom[21][36] = 8'd5;
        rom[21][37] = 8'd2;
        rom[21][38] = -8'd6;
        rom[21][39] = 8'd4;
        rom[21][40] = 8'd1;
        rom[21][41] = 8'd10;
        rom[21][42] = -8'd11;
        rom[21][43] = 8'd0;
        rom[21][44] = 8'd5;
        rom[21][45] = 8'd3;
        rom[21][46] = -8'd5;
        rom[21][47] = 8'd1;
        rom[21][48] = 8'd8;
        rom[21][49] = 8'd2;
        rom[21][50] = 8'd4;
        rom[21][51] = 8'd9;
        rom[21][52] = -8'd7;
        rom[21][53] = 8'd8;
        rom[21][54] = -8'd8;
        rom[21][55] = 8'd1;
        rom[21][56] = 8'd8;
        rom[21][57] = 8'd9;
        rom[21][58] = 8'd9;
        rom[21][59] = 8'd2;
        rom[21][60] = -8'd8;
        rom[21][61] = -8'd3;
        rom[21][62] = 8'd1;
        rom[21][63] = -8'd2;
        rom[22][0] = 8'd14;
        rom[22][1] = -8'd3;
        rom[22][2] = -8'd33;
        rom[22][3] = -8'd3;
        rom[22][4] = 8'd16;
        rom[22][5] = 8'd26;
        rom[22][6] = -8'd24;
        rom[22][7] = 8'd31;
        rom[22][8] = 8'd8;
        rom[22][9] = 8'd6;
        rom[22][10] = 8'd24;
        rom[22][11] = -8'd48;
        rom[22][12] = -8'd108;
        rom[22][13] = 8'd17;
        rom[22][14] = 8'd13;
        rom[22][15] = 8'd8;
        rom[22][16] = -8'd55;
        rom[22][17] = -8'd55;
        rom[22][18] = -8'd38;
        rom[22][19] = 8'd7;
        rom[22][20] = -8'd6;
        rom[22][21] = -8'd1;
        rom[22][22] = -8'd2;
        rom[22][23] = 8'd1;
        rom[22][24] = 8'd3;
        rom[22][25] = -8'd2;
        rom[22][26] = -8'd2;
        rom[22][27] = -8'd23;
        rom[22][28] = 8'd16;
        rom[22][29] = 8'd23;
        rom[22][30] = -8'd47;
        rom[22][31] = 8'd23;
        rom[22][32] = -8'd7;
        rom[22][33] = -8'd13;
        rom[22][34] = -8'd25;
        rom[22][35] = 8'd24;
        rom[22][36] = -8'd32;
        rom[22][37] = 8'd17;
        rom[22][38] = 8'd12;
        rom[22][39] = -8'd64;
        rom[22][40] = 8'd0;
        rom[22][41] = -8'd38;
        rom[22][42] = -8'd29;
        rom[22][43] = 8'd27;
        rom[22][44] = 8'd10;
        rom[22][45] = 8'd12;
        rom[22][46] = -8'd9;
        rom[22][47] = -8'd4;
        rom[22][48] = -8'd1;
        rom[22][49] = 8'd18;
        rom[22][50] = -8'd4;
        rom[22][51] = 8'd26;
        rom[22][52] = 8'd27;
        rom[22][53] = 8'd48;
        rom[22][54] = -8'd33;
        rom[22][55] = 8'd18;
        rom[22][56] = -8'd22;
        rom[22][57] = 8'd37;
        rom[22][58] = 8'd24;
        rom[22][59] = -8'd22;
        rom[22][60] = -8'd10;
        rom[22][61] = -8'd11;
        rom[22][62] = 8'd0;
        rom[22][63] = 8'd31;
        rom[23][0] = 8'd6;
        rom[23][1] = -8'd20;
        rom[23][2] = -8'd47;
        rom[23][3] = -8'd41;
        rom[23][4] = -8'd3;
        rom[23][5] = 8'd25;
        rom[23][6] = 8'd21;
        rom[23][7] = 8'd4;
        rom[23][8] = -8'd5;
        rom[23][9] = -8'd3;
        rom[23][10] = -8'd35;
        rom[23][11] = 8'd7;
        rom[23][12] = -8'd3;
        rom[23][13] = 8'd0;
        rom[23][14] = -8'd18;
        rom[23][15] = 8'd10;
        rom[23][16] = -8'd14;
        rom[23][17] = -8'd20;
        rom[23][18] = 8'd16;
        rom[23][19] = 8'd14;
        rom[23][20] = -8'd8;
        rom[23][21] = -8'd7;
        rom[23][22] = -8'd27;
        rom[23][23] = -8'd16;
        rom[23][24] = 8'd25;
        rom[23][25] = -8'd5;
        rom[23][26] = 8'd0;
        rom[23][27] = -8'd21;
        rom[23][28] = 8'd23;
        rom[23][29] = -8'd6;
        rom[23][30] = -8'd42;
        rom[23][31] = 8'd36;
        rom[23][32] = 8'd3;
        rom[23][33] = -8'd7;
        rom[23][34] = -8'd22;
        rom[23][35] = 8'd13;
        rom[23][36] = 8'd13;
        rom[23][37] = 8'd31;
        rom[23][38] = 8'd9;
        rom[23][39] = -8'd30;
        rom[23][40] = 8'd8;
        rom[23][41] = -8'd7;
        rom[23][42] = 8'd16;
        rom[23][43] = -8'd20;
        rom[23][44] = 8'd27;
        rom[23][45] = -8'd5;
        rom[23][46] = 8'd12;
        rom[23][47] = 8'd3;
        rom[23][48] = -8'd14;
        rom[23][49] = -8'd51;
        rom[23][50] = -8'd14;
        rom[23][51] = -8'd37;
        rom[23][52] = 8'd33;
        rom[23][53] = -8'd3;
        rom[23][54] = -8'd62;
        rom[23][55] = 8'd13;
        rom[23][56] = -8'd12;
        rom[23][57] = -8'd5;
        rom[23][58] = 8'd23;
        rom[23][59] = -8'd27;
        rom[23][60] = 8'd44;
        rom[23][61] = -8'd52;
        rom[23][62] = 8'd11;
        rom[23][63] = -8'd18;
        rom[24][0] = -8'd17;
        rom[24][1] = 8'd2;
        rom[24][2] = -8'd6;
        rom[24][3] = -8'd26;
        rom[24][4] = -8'd26;
        rom[24][5] = 8'd28;
        rom[24][6] = -8'd19;
        rom[24][7] = 8'd15;
        rom[24][8] = 8'd21;
        rom[24][9] = 8'd1;
        rom[24][10] = 8'd38;
        rom[24][11] = -8'd3;
        rom[24][12] = -8'd47;
        rom[24][13] = 8'd11;
        rom[24][14] = -8'd27;
        rom[24][15] = 8'd3;
        rom[24][16] = 8'd22;
        rom[24][17] = 8'd2;
        rom[24][18] = 8'd47;
        rom[24][19] = 8'd17;
        rom[24][20] = -8'd3;
        rom[24][21] = -8'd5;
        rom[24][22] = 8'd32;
        rom[24][23] = -8'd16;
        rom[24][24] = -8'd33;
        rom[24][25] = 8'd15;
        rom[24][26] = 8'd29;
        rom[24][27] = 8'd34;
        rom[24][28] = -8'd2;
        rom[24][29] = -8'd11;
        rom[24][30] = -8'd10;
        rom[24][31] = 8'd25;
        rom[24][32] = -8'd28;
        rom[24][33] = 8'd23;
        rom[24][34] = 8'd22;
        rom[24][35] = 8'd44;
        rom[24][36] = -8'd14;
        rom[24][37] = -8'd31;
        rom[24][38] = -8'd6;
        rom[24][39] = -8'd22;
        rom[24][40] = -8'd2;
        rom[24][41] = 8'd56;
        rom[24][42] = 8'd10;
        rom[24][43] = 8'd7;
        rom[24][44] = 8'd10;
        rom[24][45] = 8'd29;
        rom[24][46] = 8'd32;
        rom[24][47] = -8'd47;
        rom[24][48] = 8'd14;
        rom[24][49] = 8'd20;
        rom[24][50] = 8'd5;
        rom[24][51] = 8'd31;
        rom[24][52] = 8'd15;
        rom[24][53] = 8'd12;
        rom[24][54] = 8'd13;
        rom[24][55] = -8'd50;
        rom[24][56] = 8'd20;
        rom[24][57] = -8'd7;
        rom[24][58] = -8'd27;
        rom[24][59] = -8'd52;
        rom[24][60] = -8'd1;
        rom[24][61] = -8'd2;
        rom[24][62] = -8'd31;
        rom[24][63] = 8'd14;
        rom[25][0] = -8'd33;
        rom[25][1] = -8'd6;
        rom[25][2] = -8'd28;
        rom[25][3] = 8'd19;
        rom[25][4] = 8'd22;
        rom[25][5] = 8'd29;
        rom[25][6] = -8'd24;
        rom[25][7] = 8'd1;
        rom[25][8] = 8'd49;
        rom[25][9] = -8'd5;
        rom[25][10] = -8'd3;
        rom[25][11] = -8'd23;
        rom[25][12] = 8'd14;
        rom[25][13] = -8'd25;
        rom[25][14] = -8'd29;
        rom[25][15] = -8'd19;
        rom[25][16] = 8'd46;
        rom[25][17] = -8'd19;
        rom[25][18] = -8'd39;
        rom[25][19] = 8'd24;
        rom[25][20] = -8'd9;
        rom[25][21] = 8'd41;
        rom[25][22] = -8'd46;
        rom[25][23] = -8'd17;
        rom[25][24] = -8'd32;
        rom[25][25] = 8'd7;
        rom[25][26] = 8'd22;
        rom[25][27] = -8'd5;
        rom[25][28] = -8'd27;
        rom[25][29] = -8'd43;
        rom[25][30] = 8'd29;
        rom[25][31] = -8'd5;
        rom[25][32] = -8'd6;
        rom[25][33] = -8'd17;
        rom[25][34] = 8'd21;
        rom[25][35] = 8'd13;
        rom[25][36] = 8'd5;
        rom[25][37] = 8'd2;
        rom[25][38] = 8'd23;
        rom[25][39] = -8'd8;
        rom[25][40] = 8'd53;
        rom[25][41] = 8'd33;
        rom[25][42] = -8'd5;
        rom[25][43] = 8'd61;
        rom[25][44] = 8'd5;
        rom[25][45] = 8'd17;
        rom[25][46] = 8'd12;
        rom[25][47] = -8'd10;
        rom[25][48] = -8'd22;
        rom[25][49] = 8'd21;
        rom[25][50] = 8'd3;
        rom[25][51] = 8'd36;
        rom[25][52] = -8'd12;
        rom[25][53] = 8'd9;
        rom[25][54] = -8'd5;
        rom[25][55] = -8'd21;
        rom[25][56] = 8'd24;
        rom[25][57] = -8'd2;
        rom[25][58] = 8'd16;
        rom[25][59] = -8'd38;
        rom[25][60] = -8'd24;
        rom[25][61] = 8'd22;
        rom[25][62] = 8'd4;
        rom[25][63] = -8'd22;
        rom[26][0] = -8'd42;
        rom[26][1] = -8'd2;
        rom[26][2] = 8'd2;
        rom[26][3] = -8'd19;
        rom[26][4] = -8'd19;
        rom[26][5] = 8'd14;
        rom[26][6] = 8'd39;
        rom[26][7] = 8'd22;
        rom[26][8] = 8'd14;
        rom[26][9] = 8'd12;
        rom[26][10] = 8'd17;
        rom[26][11] = -8'd6;
        rom[26][12] = -8'd24;
        rom[26][13] = -8'd6;
        rom[26][14] = -8'd12;
        rom[26][15] = -8'd27;
        rom[26][16] = -8'd19;
        rom[26][17] = -8'd4;
        rom[26][18] = -8'd38;
        rom[26][19] = 8'd16;
        rom[26][20] = -8'd9;
        rom[26][21] = -8'd17;
        rom[26][22] = -8'd51;
        rom[26][23] = -8'd16;
        rom[26][24] = -8'd6;
        rom[26][25] = -8'd28;
        rom[26][26] = -8'd10;
        rom[26][27] = 8'd45;
        rom[26][28] = -8'd5;
        rom[26][29] = -8'd68;
        rom[26][30] = -8'd5;
        rom[26][31] = -8'd25;
        rom[26][32] = -8'd19;
        rom[26][33] = 8'd9;
        rom[26][34] = -8'd40;
        rom[26][35] = 8'd10;
        rom[26][36] = 8'd8;
        rom[26][37] = -8'd13;
        rom[26][38] = 8'd9;
        rom[26][39] = 8'd10;
        rom[26][40] = -8'd28;
        rom[26][41] = 8'd11;
        rom[26][42] = 8'd14;
        rom[26][43] = -8'd27;
        rom[26][44] = 8'd32;
        rom[26][45] = 8'd24;
        rom[26][46] = 8'd82;
        rom[26][47] = -8'd46;
        rom[26][48] = -8'd65;
        rom[26][49] = -8'd35;
        rom[26][50] = 8'd16;
        rom[26][51] = 8'd34;
        rom[26][52] = -8'd6;
        rom[26][53] = -8'd15;
        rom[26][54] = -8'd33;
        rom[26][55] = -8'd11;
        rom[26][56] = -8'd7;
        rom[26][57] = -8'd66;
        rom[26][58] = 8'd26;
        rom[26][59] = 8'd18;
        rom[26][60] = -8'd18;
        rom[26][61] = -8'd18;
        rom[26][62] = -8'd24;
        rom[26][63] = -8'd20;
        rom[27][0] = 8'd1;
        rom[27][1] = -8'd37;
        rom[27][2] = -8'd13;
        rom[27][3] = 8'd21;
        rom[27][4] = 8'd23;
        rom[27][5] = -8'd18;
        rom[27][6] = -8'd13;
        rom[27][7] = 8'd19;
        rom[27][8] = 8'd40;
        rom[27][9] = 8'd31;
        rom[27][10] = -8'd24;
        rom[27][11] = -8'd39;
        rom[27][12] = -8'd20;
        rom[27][13] = 8'd5;
        rom[27][14] = 8'd0;
        rom[27][15] = -8'd4;
        rom[27][16] = 8'd10;
        rom[27][17] = -8'd52;
        rom[27][18] = -8'd8;
        rom[27][19] = -8'd36;
        rom[27][20] = 8'd1;
        rom[27][21] = -8'd7;
        rom[27][22] = 8'd11;
        rom[27][23] = -8'd9;
        rom[27][24] = -8'd6;
        rom[27][25] = 8'd4;
        rom[27][26] = -8'd4;
        rom[27][27] = -8'd32;
        rom[27][28] = 8'd7;
        rom[27][29] = 8'd0;
        rom[27][30] = 8'd18;
        rom[27][31] = -8'd3;
        rom[27][32] = -8'd18;
        rom[27][33] = -8'd63;
        rom[27][34] = -8'd14;
        rom[27][35] = 8'd28;
        rom[27][36] = -8'd25;
        rom[27][37] = 8'd7;
        rom[27][38] = 8'd29;
        rom[27][39] = -8'd20;
        rom[27][40] = 8'd38;
        rom[27][41] = 8'd44;
        rom[27][42] = -8'd26;
        rom[27][43] = 8'd27;
        rom[27][44] = 8'd21;
        rom[27][45] = 8'd24;
        rom[27][46] = -8'd5;
        rom[27][47] = -8'd9;
        rom[27][48] = -8'd4;
        rom[27][49] = -8'd15;
        rom[27][50] = 8'd0;
        rom[27][51] = 8'd6;
        rom[27][52] = 8'd24;
        rom[27][53] = 8'd51;
        rom[27][54] = 8'd1;
        rom[27][55] = -8'd7;
        rom[27][56] = 8'd29;
        rom[27][57] = -8'd22;
        rom[27][58] = 8'd18;
        rom[27][59] = -8'd58;
        rom[27][60] = 8'd34;
        rom[27][61] = -8'd12;
        rom[27][62] = -8'd47;
        rom[27][63] = 8'd31;
        rom[28][0] = -8'd28;
        rom[28][1] = 8'd35;
        rom[28][2] = 8'd3;
        rom[28][3] = -8'd31;
        rom[28][4] = 8'd10;
        rom[28][5] = -8'd21;
        rom[28][6] = 8'd26;
        rom[28][7] = -8'd4;
        rom[28][8] = 8'd7;
        rom[28][9] = 8'd20;
        rom[28][10] = -8'd21;
        rom[28][11] = 8'd32;
        rom[28][12] = -8'd67;
        rom[28][13] = -8'd34;
        rom[28][14] = -8'd9;
        rom[28][15] = -8'd12;
        rom[28][16] = -8'd19;
        rom[28][17] = 8'd6;
        rom[28][18] = -8'd8;
        rom[28][19] = -8'd51;
        rom[28][20] = -8'd3;
        rom[28][21] = 8'd20;
        rom[28][22] = 8'd16;
        rom[28][23] = -8'd17;
        rom[28][24] = 8'd12;
        rom[28][25] = 8'd0;
        rom[28][26] = -8'd18;
        rom[28][27] = 8'd1;
        rom[28][28] = 8'd8;
        rom[28][29] = -8'd8;
        rom[28][30] = -8'd1;
        rom[28][31] = 8'd5;
        rom[28][32] = -8'd22;
        rom[28][33] = -8'd59;
        rom[28][34] = 8'd16;
        rom[28][35] = 8'd12;
        rom[28][36] = -8'd13;
        rom[28][37] = -8'd2;
        rom[28][38] = -8'd37;
        rom[28][39] = -8'd13;
        rom[28][40] = -8'd6;
        rom[28][41] = 8'd53;
        rom[28][42] = 8'd35;
        rom[28][43] = 8'd45;
        rom[28][44] = -8'd7;
        rom[28][45] = 8'd17;
        rom[28][46] = 8'd2;
        rom[28][47] = -8'd14;
        rom[28][48] = -8'd15;
        rom[28][49] = 8'd19;
        rom[28][50] = 8'd5;
        rom[28][51] = 8'd36;
        rom[28][52] = 8'd0;
        rom[28][53] = -8'd41;
        rom[28][54] = -8'd17;
        rom[28][55] = -8'd8;
        rom[28][56] = 8'd49;
        rom[28][57] = 8'd17;
        rom[28][58] = -8'd3;
        rom[28][59] = -8'd56;
        rom[28][60] = 8'd3;
        rom[28][61] = 8'd6;
        rom[28][62] = -8'd31;
        rom[28][63] = -8'd4;
        rom[29][0] = 8'd36;
        rom[29][1] = 8'd4;
        rom[29][2] = -8'd47;
        rom[29][3] = 8'd0;
        rom[29][4] = -8'd11;
        rom[29][5] = -8'd25;
        rom[29][6] = -8'd46;
        rom[29][7] = 8'd7;
        rom[29][8] = -8'd9;
        rom[29][9] = -8'd21;
        rom[29][10] = 8'd49;
        rom[29][11] = 8'd22;
        rom[29][12] = -8'd31;
        rom[29][13] = 8'd8;
        rom[29][14] = -8'd17;
        rom[29][15] = 8'd24;
        rom[29][16] = -8'd10;
        rom[29][17] = 8'd28;
        rom[29][18] = 8'd2;
        rom[29][19] = 8'd11;
        rom[29][20] = -8'd3;
        rom[29][21] = 8'd6;
        rom[29][22] = 8'd14;
        rom[29][23] = -8'd108;
        rom[29][24] = -8'd42;
        rom[29][25] = 8'd9;
        rom[29][26] = -8'd7;
        rom[29][27] = -8'd52;
        rom[29][28] = 8'd34;
        rom[29][29] = -8'd12;
        rom[29][30] = -8'd2;
        rom[29][31] = 8'd15;
        rom[29][32] = -8'd19;
        rom[29][33] = -8'd65;
        rom[29][34] = -8'd13;
        rom[29][35] = 8'd22;
        rom[29][36] = -8'd7;
        rom[29][37] = 8'd0;
        rom[29][38] = -8'd10;
        rom[29][39] = 8'd7;
        rom[29][40] = -8'd26;
        rom[29][41] = 8'd17;
        rom[29][42] = -8'd28;
        rom[29][43] = -8'd34;
        rom[29][44] = -8'd26;
        rom[29][45] = -8'd6;
        rom[29][46] = -8'd1;
        rom[29][47] = 8'd44;
        rom[29][48] = 8'd4;
        rom[29][49] = -8'd9;
        rom[29][50] = -8'd23;
        rom[29][51] = 8'd29;
        rom[29][52] = -8'd25;
        rom[29][53] = -8'd52;
        rom[29][54] = 8'd6;
        rom[29][55] = -8'd21;
        rom[29][56] = 8'd27;
        rom[29][57] = -8'd8;
        rom[29][58] = -8'd73;
        rom[29][59] = -8'd51;
        rom[29][60] = -8'd5;
        rom[29][61] = -8'd7;
        rom[29][62] = -8'd20;
        rom[29][63] = 8'd33;
        rom[30][0] = -8'd4;
        rom[30][1] = 8'd3;
        rom[30][2] = 8'd28;
        rom[30][3] = -8'd16;
        rom[30][4] = 8'd25;
        rom[30][5] = -8'd37;
        rom[30][6] = 8'd5;
        rom[30][7] = -8'd14;
        rom[30][8] = 8'd20;
        rom[30][9] = 8'd32;
        rom[30][10] = -8'd16;
        rom[30][11] = -8'd14;
        rom[30][12] = 8'd21;
        rom[30][13] = 8'd1;
        rom[30][14] = -8'd8;
        rom[30][15] = 8'd4;
        rom[30][16] = 8'd0;
        rom[30][17] = 8'd3;
        rom[30][18] = -8'd61;
        rom[30][19] = -8'd14;
        rom[30][20] = -8'd7;
        rom[30][21] = -8'd1;
        rom[30][22] = -8'd19;
        rom[30][23] = -8'd20;
        rom[30][24] = 8'd5;
        rom[30][25] = -8'd82;
        rom[30][26] = -8'd32;
        rom[30][27] = 8'd3;
        rom[30][28] = -8'd87;
        rom[30][29] = 8'd24;
        rom[30][30] = 8'd14;
        rom[30][31] = 8'd8;
        rom[30][32] = 8'd20;
        rom[30][33] = 8'd12;
        rom[30][34] = 8'd5;
        rom[30][35] = 8'd6;
        rom[30][36] = 8'd22;
        rom[30][37] = -8'd8;
        rom[30][38] = 8'd21;
        rom[30][39] = 8'd7;
        rom[30][40] = 8'd8;
        rom[30][41] = 8'd28;
        rom[30][42] = -8'd19;
        rom[30][43] = -8'd18;
        rom[30][44] = -8'd66;
        rom[30][45] = -8'd12;
        rom[30][46] = -8'd5;
        rom[30][47] = 8'd29;
        rom[30][48] = -8'd29;
        rom[30][49] = 8'd21;
        rom[30][50] = -8'd18;
        rom[30][51] = 8'd9;
        rom[30][52] = -8'd43;
        rom[30][53] = 8'd29;
        rom[30][54] = -8'd40;
        rom[30][55] = 8'd20;
        rom[30][56] = 8'd46;
        rom[30][57] = 8'd11;
        rom[30][58] = -8'd59;
        rom[30][59] = -8'd15;
        rom[30][60] = -8'd6;
        rom[30][61] = -8'd5;
        rom[30][62] = -8'd56;
        rom[30][63] = -8'd18;
        rom[31][0] = 8'd3;
        rom[31][1] = -8'd126;
        rom[31][2] = 8'd14;
        rom[31][3] = -8'd41;
        rom[31][4] = 8'd5;
        rom[31][5] = -8'd7;
        rom[31][6] = 8'd35;
        rom[31][7] = 8'd43;
        rom[31][8] = 8'd3;
        rom[31][9] = -8'd6;
        rom[31][10] = -8'd15;
        rom[31][11] = -8'd76;
        rom[31][12] = 8'd3;
        rom[31][13] = -8'd37;
        rom[31][14] = 8'd19;
        rom[31][15] = 8'd11;
        rom[31][16] = 8'd19;
        rom[31][17] = -8'd4;
        rom[31][18] = 8'd4;
        rom[31][19] = 8'd18;
        rom[31][20] = -8'd9;
        rom[31][21] = -8'd45;
        rom[31][22] = 8'd7;
        rom[31][23] = -8'd23;
        rom[31][24] = -8'd22;
        rom[31][25] = 8'd45;
        rom[31][26] = -8'd33;
        rom[31][27] = -8'd17;
        rom[31][28] = 8'd19;
        rom[31][29] = -8'd3;
        rom[31][30] = -8'd13;
        rom[31][31] = -8'd28;
        rom[31][32] = -8'd47;
        rom[31][33] = 8'd15;
        rom[31][34] = 8'd41;
        rom[31][35] = -8'd2;
        rom[31][36] = 8'd10;
        rom[31][37] = -8'd43;
        rom[31][38] = -8'd15;
        rom[31][39] = 8'd26;
        rom[31][40] = -8'd6;
        rom[31][41] = -8'd40;
        rom[31][42] = 8'd21;
        rom[31][43] = 8'd10;
        rom[31][44] = 8'd6;
        rom[31][45] = -8'd39;
        rom[31][46] = 8'd2;
        rom[31][47] = -8'd14;
        rom[31][48] = -8'd12;
        rom[31][49] = -8'd3;
        rom[31][50] = 8'd20;
        rom[31][51] = 8'd3;
        rom[31][52] = 8'd40;
        rom[31][53] = 8'd21;
        rom[31][54] = 8'd25;
        rom[31][55] = -8'd40;
        rom[31][56] = -8'd38;
        rom[31][57] = -8'd19;
        rom[31][58] = 8'd10;
        rom[31][59] = 8'd11;
        rom[31][60] = 8'd10;
        rom[31][61] = -8'd2;
        rom[31][62] = -8'd26;
        rom[31][63] = 8'd6;
        rom[32][0] = -8'd11;
        rom[32][1] = 8'd24;
        rom[32][2] = 8'd2;
        rom[32][3] = -8'd32;
        rom[32][4] = 8'd7;
        rom[32][5] = 8'd25;
        rom[32][6] = -8'd10;
        rom[32][7] = -8'd26;
        rom[32][8] = -8'd5;
        rom[32][9] = -8'd21;
        rom[32][10] = -8'd29;
        rom[32][11] = -8'd38;
        rom[32][12] = -8'd1;
        rom[32][13] = 8'd10;
        rom[32][14] = 8'd34;
        rom[32][15] = -8'd10;
        rom[32][16] = -8'd14;
        rom[32][17] = -8'd15;
        rom[32][18] = -8'd14;
        rom[32][19] = 8'd2;
        rom[32][20] = 8'd4;
        rom[32][21] = 8'd24;
        rom[32][22] = 8'd13;
        rom[32][23] = 8'd4;
        rom[32][24] = -8'd44;
        rom[32][25] = -8'd18;
        rom[32][26] = -8'd65;
        rom[32][27] = -8'd30;
        rom[32][28] = -8'd24;
        rom[32][29] = -8'd43;
        rom[32][30] = -8'd15;
        rom[32][31] = -8'd26;
        rom[32][32] = -8'd3;
        rom[32][33] = 8'd41;
        rom[32][34] = -8'd67;
        rom[32][35] = -8'd11;
        rom[32][36] = -8'd3;
        rom[32][37] = 8'd4;
        rom[32][38] = -8'd26;
        rom[32][39] = 8'd0;
        rom[32][40] = 8'd11;
        rom[32][41] = -8'd25;
        rom[32][42] = 8'd19;
        rom[32][43] = -8'd15;
        rom[32][44] = -8'd11;
        rom[32][45] = 8'd8;
        rom[32][46] = 8'd26;
        rom[32][47] = 8'd0;
        rom[32][48] = 8'd12;
        rom[32][49] = 8'd24;
        rom[32][50] = -8'd8;
        rom[32][51] = -8'd9;
        rom[32][52] = 8'd30;
        rom[32][53] = -8'd25;
        rom[32][54] = -8'd13;
        rom[32][55] = -8'd51;
        rom[32][56] = -8'd6;
        rom[32][57] = -8'd40;
        rom[32][58] = -8'd4;
        rom[32][59] = -8'd2;
        rom[32][60] = -8'd50;
        rom[32][61] = -8'd26;
        rom[32][62] = -8'd39;
        rom[32][63] = -8'd29;
        rom[33][0] = 8'd20;
        rom[33][1] = 8'd66;
        rom[33][2] = 8'd7;
        rom[33][3] = 8'd36;
        rom[33][4] = -8'd39;
        rom[33][5] = 8'd12;
        rom[33][6] = 8'd46;
        rom[33][7] = 8'd29;
        rom[33][8] = 8'd36;
        rom[33][9] = -8'd2;
        rom[33][10] = 8'd32;
        rom[33][11] = 8'd25;
        rom[33][12] = 8'd30;
        rom[33][13] = -8'd60;
        rom[33][14] = -8'd42;
        rom[33][15] = 8'd19;
        rom[33][16] = 8'd5;
        rom[33][17] = 8'd11;
        rom[33][18] = 8'd30;
        rom[33][19] = -8'd16;
        rom[33][20] = -8'd7;
        rom[33][21] = -8'd10;
        rom[33][22] = -8'd32;
        rom[33][23] = 8'd10;
        rom[33][24] = -8'd30;
        rom[33][25] = 8'd24;
        rom[33][26] = -8'd37;
        rom[33][27] = 8'd8;
        rom[33][28] = -8'd16;
        rom[33][29] = -8'd20;
        rom[33][30] = 8'd1;
        rom[33][31] = -8'd15;
        rom[33][32] = -8'd26;
        rom[33][33] = -8'd55;
        rom[33][34] = -8'd62;
        rom[33][35] = -8'd33;
        rom[33][36] = 8'd58;
        rom[33][37] = -8'd3;
        rom[33][38] = 8'd48;
        rom[33][39] = 8'd21;
        rom[33][40] = -8'd3;
        rom[33][41] = -8'd27;
        rom[33][42] = -8'd4;
        rom[33][43] = 8'd8;
        rom[33][44] = -8'd41;
        rom[33][45] = 8'd40;
        rom[33][46] = -8'd20;
        rom[33][47] = -8'd24;
        rom[33][48] = -8'd7;
        rom[33][49] = -8'd6;
        rom[33][50] = -8'd38;
        rom[33][51] = 8'd12;
        rom[33][52] = -8'd75;
        rom[33][53] = -8'd45;
        rom[33][54] = 8'd9;
        rom[33][55] = 8'd33;
        rom[33][56] = -8'd70;
        rom[33][57] = -8'd4;
        rom[33][58] = 8'd20;
        rom[33][59] = 8'd38;
        rom[33][60] = 8'd70;
        rom[33][61] = 8'd20;
        rom[33][62] = 8'd3;
        rom[33][63] = -8'd51;
        rom[34][0] = 8'd17;
        rom[34][1] = 8'd32;
        rom[34][2] = 8'd0;
        rom[34][3] = 8'd42;
        rom[34][4] = -8'd5;
        rom[34][5] = -8'd5;
        rom[34][6] = 8'd13;
        rom[34][7] = 8'd1;
        rom[34][8] = 8'd44;
        rom[34][9] = 8'd28;
        rom[34][10] = 8'd26;
        rom[34][11] = 8'd47;
        rom[34][12] = -8'd32;
        rom[34][13] = -8'd23;
        rom[34][14] = 8'd45;
        rom[34][15] = -8'd12;
        rom[34][16] = -8'd14;
        rom[34][17] = -8'd14;
        rom[34][18] = 8'd17;
        rom[34][19] = -8'd15;
        rom[34][20] = -8'd9;
        rom[34][21] = -8'd8;
        rom[34][22] = 8'd42;
        rom[34][23] = 8'd0;
        rom[34][24] = 8'd36;
        rom[34][25] = 8'd5;
        rom[34][26] = -8'd13;
        rom[34][27] = -8'd128;
        rom[34][28] = -8'd48;
        rom[34][29] = -8'd4;
        rom[34][30] = 8'd7;
        rom[34][31] = 8'd0;
        rom[34][32] = -8'd3;
        rom[34][33] = -8'd49;
        rom[34][34] = 8'd6;
        rom[34][35] = 8'd5;
        rom[34][36] = 8'd25;
        rom[34][37] = -8'd22;
        rom[34][38] = 8'd17;
        rom[34][39] = 8'd39;
        rom[34][40] = 8'd2;
        rom[34][41] = -8'd16;
        rom[34][42] = 8'd26;
        rom[34][43] = -8'd76;
        rom[34][44] = -8'd48;
        rom[34][45] = -8'd7;
        rom[34][46] = 8'd21;
        rom[34][47] = -8'd40;
        rom[34][48] = -8'd9;
        rom[34][49] = 8'd50;
        rom[34][50] = -8'd27;
        rom[34][51] = 8'd26;
        rom[34][52] = -8'd2;
        rom[34][53] = -8'd11;
        rom[34][54] = -8'd11;
        rom[34][55] = -8'd6;
        rom[34][56] = -8'd19;
        rom[34][57] = -8'd12;
        rom[34][58] = -8'd128;
        rom[34][59] = -8'd2;
        rom[34][60] = -8'd29;
        rom[34][61] = 8'd49;
        rom[34][62] = -8'd2;
        rom[34][63] = -8'd2;
        rom[35][0] = 8'd34;
        rom[35][1] = 8'd23;
        rom[35][2] = 8'd29;
        rom[35][3] = -8'd54;
        rom[35][4] = -8'd27;
        rom[35][5] = -8'd55;
        rom[35][6] = -8'd13;
        rom[35][7] = -8'd20;
        rom[35][8] = 8'd11;
        rom[35][9] = 8'd3;
        rom[35][10] = -8'd46;
        rom[35][11] = 8'd16;
        rom[35][12] = 8'd33;
        rom[35][13] = -8'd39;
        rom[35][14] = 8'd8;
        rom[35][15] = 8'd11;
        rom[35][16] = 8'd48;
        rom[35][17] = -8'd41;
        rom[35][18] = -8'd34;
        rom[35][19] = -8'd63;
        rom[35][20] = -8'd13;
        rom[35][21] = -8'd36;
        rom[35][22] = 8'd3;
        rom[35][23] = 8'd23;
        rom[35][24] = -8'd23;
        rom[35][25] = 8'd12;
        rom[35][26] = -8'd55;
        rom[35][27] = 8'd5;
        rom[35][28] = -8'd18;
        rom[35][29] = 8'd32;
        rom[35][30] = -8'd63;
        rom[35][31] = 8'd11;
        rom[35][32] = 8'd6;
        rom[35][33] = -8'd48;
        rom[35][34] = 8'd3;
        rom[35][35] = 8'd34;
        rom[35][36] = 8'd4;
        rom[35][37] = 8'd15;
        rom[35][38] = 8'd4;
        rom[35][39] = -8'd25;
        rom[35][40] = -8'd44;
        rom[35][41] = -8'd50;
        rom[35][42] = -8'd60;
        rom[35][43] = 8'd13;
        rom[35][44] = -8'd10;
        rom[35][45] = -8'd9;
        rom[35][46] = 8'd15;
        rom[35][47] = 8'd3;
        rom[35][48] = -8'd20;
        rom[35][49] = 8'd2;
        rom[35][50] = 8'd27;
        rom[35][51] = 8'd24;
        rom[35][52] = -8'd16;
        rom[35][53] = -8'd15;
        rom[35][54] = 8'd17;
        rom[35][55] = -8'd23;
        rom[35][56] = -8'd4;
        rom[35][57] = -8'd4;
        rom[35][58] = 8'd3;
        rom[35][59] = 8'd15;
        rom[35][60] = -8'd3;
        rom[35][61] = 8'd2;
        rom[35][62] = -8'd26;
        rom[35][63] = 8'd4;
        rom[36][0] = -8'd40;
        rom[36][1] = -8'd32;
        rom[36][2] = 8'd9;
        rom[36][3] = 8'd1;
        rom[36][4] = 8'd12;
        rom[36][5] = -8'd15;
        rom[36][6] = 8'd2;
        rom[36][7] = 8'd13;
        rom[36][8] = 8'd30;
        rom[36][9] = -8'd10;
        rom[36][10] = -8'd11;
        rom[36][11] = 8'd6;
        rom[36][12] = -8'd83;
        rom[36][13] = -8'd4;
        rom[36][14] = -8'd12;
        rom[36][15] = 8'd39;
        rom[36][16] = -8'd64;
        rom[36][17] = 8'd0;
        rom[36][18] = 8'd1;
        rom[36][19] = 8'd10;
        rom[36][20] = -8'd9;
        rom[36][21] = 8'd6;
        rom[36][22] = 8'd16;
        rom[36][23] = -8'd24;
        rom[36][24] = -8'd13;
        rom[36][25] = 8'd9;
        rom[36][26] = -8'd23;
        rom[36][27] = 8'd9;
        rom[36][28] = -8'd14;
        rom[36][29] = -8'd2;
        rom[36][30] = -8'd14;
        rom[36][31] = 8'd11;
        rom[36][32] = -8'd52;
        rom[36][33] = -8'd29;
        rom[36][34] = -8'd14;
        rom[36][35] = 8'd6;
        rom[36][36] = -8'd4;
        rom[36][37] = 8'd27;
        rom[36][38] = -8'd8;
        rom[36][39] = -8'd6;
        rom[36][40] = -8'd8;
        rom[36][41] = -8'd49;
        rom[36][42] = 8'd9;
        rom[36][43] = 8'd24;
        rom[36][44] = -8'd11;
        rom[36][45] = 8'd8;
        rom[36][46] = 8'd5;
        rom[36][47] = 8'd0;
        rom[36][48] = 8'd5;
        rom[36][49] = 8'd7;
        rom[36][50] = 8'd16;
        rom[36][51] = -8'd27;
        rom[36][52] = -8'd12;
        rom[36][53] = 8'd22;
        rom[36][54] = 8'd17;
        rom[36][55] = 8'd36;
        rom[36][56] = -8'd43;
        rom[36][57] = -8'd41;
        rom[36][58] = 8'd28;
        rom[36][59] = 8'd17;
        rom[36][60] = 8'd11;
        rom[36][61] = -8'd20;
        rom[36][62] = 8'd0;
        rom[36][63] = -8'd7;
        rom[37][0] = -8'd12;
        rom[37][1] = -8'd45;
        rom[37][2] = -8'd20;
        rom[37][3] = -8'd20;
        rom[37][4] = 8'd6;
        rom[37][5] = -8'd2;
        rom[37][6] = -8'd14;
        rom[37][7] = 8'd18;
        rom[37][8] = 8'd16;
        rom[37][9] = 8'd15;
        rom[37][10] = -8'd49;
        rom[37][11] = -8'd22;
        rom[37][12] = -8'd5;
        rom[37][13] = -8'd30;
        rom[37][14] = 8'd23;
        rom[37][15] = 8'd24;
        rom[37][16] = -8'd76;
        rom[37][17] = 8'd15;
        rom[37][18] = -8'd7;
        rom[37][19] = -8'd8;
        rom[37][20] = -8'd6;
        rom[37][21] = -8'd8;
        rom[37][22] = 8'd17;
        rom[37][23] = -8'd44;
        rom[37][24] = 8'd13;
        rom[37][25] = 8'd22;
        rom[37][26] = -8'd4;
        rom[37][27] = 8'd27;
        rom[37][28] = -8'd20;
        rom[37][29] = -8'd5;
        rom[37][30] = 8'd1;
        rom[37][31] = -8'd24;
        rom[37][32] = -8'd22;
        rom[37][33] = -8'd41;
        rom[37][34] = -8'd30;
        rom[37][35] = 8'd14;
        rom[37][36] = -8'd19;
        rom[37][37] = 8'd18;
        rom[37][38] = -8'd104;
        rom[37][39] = -8'd25;
        rom[37][40] = 8'd2;
        rom[37][41] = 8'd23;
        rom[37][42] = -8'd30;
        rom[37][43] = 8'd2;
        rom[37][44] = -8'd51;
        rom[37][45] = 8'd40;
        rom[37][46] = -8'd42;
        rom[37][47] = 8'd5;
        rom[37][48] = -8'd13;
        rom[37][49] = -8'd1;
        rom[37][50] = 8'd16;
        rom[37][51] = -8'd11;
        rom[37][52] = -8'd10;
        rom[37][53] = 8'd22;
        rom[37][54] = 8'd2;
        rom[37][55] = 8'd9;
        rom[37][56] = -8'd2;
        rom[37][57] = -8'd6;
        rom[37][58] = -8'd15;
        rom[37][59] = -8'd15;
        rom[37][60] = 8'd1;
        rom[37][61] = 8'd7;
        rom[37][62] = -8'd23;
        rom[37][63] = -8'd25;
        rom[38][0] = -8'd43;
        rom[38][1] = 8'd36;
        rom[38][2] = 8'd51;
        rom[38][3] = -8'd7;
        rom[38][4] = -8'd22;
        rom[38][5] = -8'd9;
        rom[38][6] = -8'd35;
        rom[38][7] = -8'd14;
        rom[38][8] = -8'd45;
        rom[38][9] = 8'd31;
        rom[38][10] = -8'd28;
        rom[38][11] = -8'd43;
        rom[38][12] = 8'd19;
        rom[38][13] = -8'd24;
        rom[38][14] = -8'd2;
        rom[38][15] = -8'd35;
        rom[38][16] = 8'd32;
        rom[38][17] = -8'd1;
        rom[38][18] = 8'd4;
        rom[38][19] = -8'd22;
        rom[38][20] = -8'd2;
        rom[38][21] = -8'd40;
        rom[38][22] = -8'd98;
        rom[38][23] = -8'd51;
        rom[38][24] = -8'd34;
        rom[38][25] = 8'd11;
        rom[38][26] = 8'd23;
        rom[38][27] = -8'd71;
        rom[38][28] = 8'd31;
        rom[38][29] = 8'd8;
        rom[38][30] = 8'd40;
        rom[38][31] = 8'd40;
        rom[38][32] = 8'd9;
        rom[38][33] = -8'd96;
        rom[38][34] = 8'd20;
        rom[38][35] = 8'd20;
        rom[38][36] = -8'd18;
        rom[38][37] = 8'd7;
        rom[38][38] = -8'd31;
        rom[38][39] = -8'd33;
        rom[38][40] = -8'd16;
        rom[38][41] = -8'd28;
        rom[38][42] = 8'd30;
        rom[38][43] = 8'd47;
        rom[38][44] = 8'd20;
        rom[38][45] = -8'd71;
        rom[38][46] = -8'd29;
        rom[38][47] = 8'd24;
        rom[38][48] = 8'd27;
        rom[38][49] = -8'd29;
        rom[38][50] = -8'd54;
        rom[38][51] = 8'd10;
        rom[38][52] = 8'd7;
        rom[38][53] = 8'd8;
        rom[38][54] = 8'd44;
        rom[38][55] = -8'd86;
        rom[38][56] = 8'd1;
        rom[38][57] = 8'd32;
        rom[38][58] = -8'd71;
        rom[38][59] = -8'd27;
        rom[38][60] = 8'd9;
        rom[38][61] = -8'd41;
        rom[38][62] = 8'd36;
        rom[38][63] = -8'd36;
        rom[39][0] = -8'd13;
        rom[39][1] = 8'd24;
        rom[39][2] = -8'd8;
        rom[39][3] = 8'd27;
        rom[39][4] = -8'd13;
        rom[39][5] = 8'd19;
        rom[39][6] = -8'd18;
        rom[39][7] = 8'd2;
        rom[39][8] = 8'd18;
        rom[39][9] = -8'd21;
        rom[39][10] = 8'd6;
        rom[39][11] = 8'd0;
        rom[39][12] = 8'd12;
        rom[39][13] = 8'd14;
        rom[39][14] = 8'd10;
        rom[39][15] = -8'd11;
        rom[39][16] = -8'd2;
        rom[39][17] = 8'd6;
        rom[39][18] = 8'd25;
        rom[39][19] = 8'd24;
        rom[39][20] = -8'd3;
        rom[39][21] = -8'd22;
        rom[39][22] = -8'd32;
        rom[39][23] = -8'd42;
        rom[39][24] = -8'd10;
        rom[39][25] = -8'd35;
        rom[39][26] = 8'd4;
        rom[39][27] = -8'd28;
        rom[39][28] = -8'd5;
        rom[39][29] = -8'd4;
        rom[39][30] = 8'd13;
        rom[39][31] = -8'd22;
        rom[39][32] = -8'd9;
        rom[39][33] = -8'd70;
        rom[39][34] = -8'd4;
        rom[39][35] = 8'd28;
        rom[39][36] = -8'd1;
        rom[39][37] = -8'd20;
        rom[39][38] = -8'd29;
        rom[39][39] = 8'd4;
        rom[39][40] = 8'd1;
        rom[39][41] = -8'd5;
        rom[39][42] = 8'd31;
        rom[39][43] = 8'd0;
        rom[39][44] = -8'd11;
        rom[39][45] = -8'd2;
        rom[39][46] = 8'd14;
        rom[39][47] = -8'd37;
        rom[39][48] = -8'd9;
        rom[39][49] = 8'd26;
        rom[39][50] = -8'd19;
        rom[39][51] = -8'd21;
        rom[39][52] = -8'd10;
        rom[39][53] = 8'd5;
        rom[39][54] = -8'd7;
        rom[39][55] = -8'd44;
        rom[39][56] = -8'd2;
        rom[39][57] = -8'd30;
        rom[39][58] = -8'd26;
        rom[39][59] = 8'd4;
        rom[39][60] = 8'd8;
        rom[39][61] = -8'd28;
        rom[39][62] = 8'd31;
        rom[39][63] = -8'd12;
        rom[40][0] = -8'd23;
        rom[40][1] = -8'd54;
        rom[40][2] = -8'd35;
        rom[40][3] = -8'd9;
        rom[40][4] = -8'd7;
        rom[40][5] = -8'd2;
        rom[40][6] = 8'd12;
        rom[40][7] = 8'd14;
        rom[40][8] = -8'd2;
        rom[40][9] = -8'd65;
        rom[40][10] = -8'd109;
        rom[40][11] = 8'd2;
        rom[40][12] = -8'd7;
        rom[40][13] = -8'd8;
        rom[40][14] = -8'd26;
        rom[40][15] = -8'd38;
        rom[40][16] = -8'd5;
        rom[40][17] = -8'd27;
        rom[40][18] = -8'd16;
        rom[40][19] = 8'd17;
        rom[40][20] = -8'd5;
        rom[40][21] = -8'd28;
        rom[40][22] = -8'd2;
        rom[40][23] = 8'd25;
        rom[40][24] = 8'd37;
        rom[40][25] = -8'd44;
        rom[40][26] = -8'd21;
        rom[40][27] = -8'd13;
        rom[40][28] = -8'd20;
        rom[40][29] = -8'd60;
        rom[40][30] = -8'd5;
        rom[40][31] = 8'd58;
        rom[40][32] = 8'd19;
        rom[40][33] = -8'd9;
        rom[40][34] = 8'd40;
        rom[40][35] = 8'd17;
        rom[40][36] = -8'd10;
        rom[40][37] = -8'd32;
        rom[40][38] = 8'd29;
        rom[40][39] = -8'd2;
        rom[40][40] = 8'd24;
        rom[40][41] = 8'd29;
        rom[40][42] = 8'd41;
        rom[40][43] = 8'd17;
        rom[40][44] = 8'd9;
        rom[40][45] = 8'd1;
        rom[40][46] = 8'd24;
        rom[40][47] = 8'd26;
        rom[40][48] = 8'd38;
        rom[40][49] = -8'd24;
        rom[40][50] = -8'd12;
        rom[40][51] = -8'd4;
        rom[40][52] = -8'd30;
        rom[40][53] = -8'd17;
        rom[40][54] = 8'd31;
        rom[40][55] = 8'd1;
        rom[40][56] = -8'd6;
        rom[40][57] = 8'd2;
        rom[40][58] = 8'd41;
        rom[40][59] = 8'd8;
        rom[40][60] = -8'd43;
        rom[40][61] = -8'd40;
        rom[40][62] = 8'd54;
        rom[40][63] = 8'd12;
        rom[41][0] = -8'd6;
        rom[41][1] = -8'd19;
        rom[41][2] = 8'd15;
        rom[41][3] = 8'd35;
        rom[41][4] = 8'd40;
        rom[41][5] = 8'd25;
        rom[41][6] = 8'd6;
        rom[41][7] = -8'd11;
        rom[41][8] = 8'd8;
        rom[41][9] = 8'd19;
        rom[41][10] = -8'd3;
        rom[41][11] = -8'd17;
        rom[41][12] = -8'd21;
        rom[41][13] = 8'd26;
        rom[41][14] = -8'd12;
        rom[41][15] = -8'd25;
        rom[41][16] = -8'd40;
        rom[41][17] = -8'd76;
        rom[41][18] = -8'd52;
        rom[41][19] = -8'd21;
        rom[41][20] = 8'd5;
        rom[41][21] = -8'd45;
        rom[41][22] = -8'd32;
        rom[41][23] = 8'd17;
        rom[41][24] = 8'd43;
        rom[41][25] = -8'd31;
        rom[41][26] = -8'd21;
        rom[41][27] = -8'd22;
        rom[41][28] = 8'd23;
        rom[41][29] = -8'd8;
        rom[41][30] = 8'd28;
        rom[41][31] = 8'd19;
        rom[41][32] = -8'd34;
        rom[41][33] = -8'd35;
        rom[41][34] = 8'd7;
        rom[41][35] = 8'd1;
        rom[41][36] = -8'd14;
        rom[41][37] = -8'd17;
        rom[41][38] = -8'd26;
        rom[41][39] = 8'd3;
        rom[41][40] = 8'd5;
        rom[41][41] = -8'd35;
        rom[41][42] = 8'd29;
        rom[41][43] = 8'd10;
        rom[41][44] = -8'd9;
        rom[41][45] = -8'd11;
        rom[41][46] = 8'd10;
        rom[41][47] = -8'd22;
        rom[41][48] = 8'd23;
        rom[41][49] = -8'd7;
        rom[41][50] = 8'd10;
        rom[41][51] = 8'd19;
        rom[41][52] = 8'd1;
        rom[41][53] = -8'd3;
        rom[41][54] = -8'd32;
        rom[41][55] = -8'd4;
        rom[41][56] = -8'd17;
        rom[41][57] = 8'd9;
        rom[41][58] = 8'd16;
        rom[41][59] = 8'd7;
        rom[41][60] = 8'd22;
        rom[41][61] = -8'd9;
        rom[41][62] = -8'd2;
        rom[41][63] = 8'd17;
        rom[42][0] = -8'd4;
        rom[42][1] = -8'd5;
        rom[42][2] = 8'd27;
        rom[42][3] = -8'd31;
        rom[42][4] = -8'd40;
        rom[42][5] = 8'd13;
        rom[42][6] = 8'd10;
        rom[42][7] = 8'd24;
        rom[42][8] = 8'd25;
        rom[42][9] = 8'd11;
        rom[42][10] = 8'd27;
        rom[42][11] = 8'd3;
        rom[42][12] = -8'd6;
        rom[42][13] = 8'd12;
        rom[42][14] = -8'd6;
        rom[42][15] = -8'd28;
        rom[42][16] = 8'd8;
        rom[42][17] = -8'd6;
        rom[42][18] = 8'd2;
        rom[42][19] = -8'd12;
        rom[42][20] = -8'd2;
        rom[42][21] = -8'd11;
        rom[42][22] = -8'd15;
        rom[42][23] = 8'd21;
        rom[42][24] = -8'd34;
        rom[42][25] = 8'd1;
        rom[42][26] = 8'd31;
        rom[42][27] = 8'd8;
        rom[42][28] = 8'd10;
        rom[42][29] = -8'd83;
        rom[42][30] = 8'd14;
        rom[42][31] = -8'd98;
        rom[42][32] = -8'd26;
        rom[42][33] = 8'd2;
        rom[42][34] = 8'd11;
        rom[42][35] = 8'd6;
        rom[42][36] = -8'd18;
        rom[42][37] = -8'd25;
        rom[42][38] = 8'd16;
        rom[42][39] = 8'd28;
        rom[42][40] = -8'd45;
        rom[42][41] = 8'd7;
        rom[42][42] = 8'd27;
        rom[42][43] = -8'd18;
        rom[42][44] = 8'd4;
        rom[42][45] = -8'd6;
        rom[42][46] = 8'd20;
        rom[42][47] = -8'd8;
        rom[42][48] = 8'd7;
        rom[42][49] = -8'd63;
        rom[42][50] = 8'd27;
        rom[42][51] = 8'd25;
        rom[42][52] = -8'd7;
        rom[42][53] = -8'd1;
        rom[42][54] = 8'd8;
        rom[42][55] = 8'd11;
        rom[42][56] = 8'd2;
        rom[42][57] = 8'd21;
        rom[42][58] = -8'd5;
        rom[42][59] = 8'd33;
        rom[42][60] = -8'd10;
        rom[42][61] = -8'd8;
        rom[42][62] = -8'd33;
        rom[42][63] = -8'd12;
        rom[43][0] = -8'd12;
        rom[43][1] = -8'd33;
        rom[43][2] = 8'd31;
        rom[43][3] = 8'd7;
        rom[43][4] = 8'd6;
        rom[43][5] = 8'd8;
        rom[43][6] = -8'd20;
        rom[43][7] = -8'd5;
        rom[43][8] = 8'd14;
        rom[43][9] = 8'd26;
        rom[43][10] = -8'd18;
        rom[43][11] = 8'd1;
        rom[43][12] = -8'd32;
        rom[43][13] = -8'd5;
        rom[43][14] = 8'd6;
        rom[43][15] = -8'd6;
        rom[43][16] = -8'd80;
        rom[43][17] = -8'd1;
        rom[43][18] = 8'd31;
        rom[43][19] = -8'd20;
        rom[43][20] = -8'd9;
        rom[43][21] = 8'd11;
        rom[43][22] = -8'd39;
        rom[43][23] = -8'd33;
        rom[43][24] = 8'd2;
        rom[43][25] = 8'd34;
        rom[43][26] = 8'd16;
        rom[43][27] = -8'd4;
        rom[43][28] = 8'd43;
        rom[43][29] = 8'd9;
        rom[43][30] = -8'd31;
        rom[43][31] = 8'd1;
        rom[43][32] = -8'd42;
        rom[43][33] = -8'd65;
        rom[43][34] = 8'd12;
        rom[43][35] = 8'd34;
        rom[43][36] = 8'd27;
        rom[43][37] = -8'd24;
        rom[43][38] = 8'd4;
        rom[43][39] = -8'd16;
        rom[43][40] = -8'd24;
        rom[43][41] = -8'd16;
        rom[43][42] = 8'd18;
        rom[43][43] = 8'd13;
        rom[43][44] = -8'd39;
        rom[43][45] = -8'd4;
        rom[43][46] = 8'd0;
        rom[43][47] = -8'd9;
        rom[43][48] = 8'd8;
        rom[43][49] = 8'd8;
        rom[43][50] = -8'd15;
        rom[43][51] = -8'd12;
        rom[43][52] = 8'd9;
        rom[43][53] = 8'd29;
        rom[43][54] = -8'd1;
        rom[43][55] = 8'd28;
        rom[43][56] = -8'd23;
        rom[43][57] = -8'd30;
        rom[43][58] = 8'd8;
        rom[43][59] = 8'd15;
        rom[43][60] = 8'd1;
        rom[43][61] = 8'd16;
        rom[43][62] = 8'd6;
        rom[43][63] = 8'd17;
        rom[44][0] = -8'd35;
        rom[44][1] = -8'd14;
        rom[44][2] = -8'd15;
        rom[44][3] = -8'd17;
        rom[44][4] = 8'd24;
        rom[44][5] = -8'd14;
        rom[44][6] = 8'd17;
        rom[44][7] = -8'd54;
        rom[44][8] = 8'd9;
        rom[44][9] = 8'd16;
        rom[44][10] = -8'd6;
        rom[44][11] = -8'd12;
        rom[44][12] = 8'd29;
        rom[44][13] = -8'd16;
        rom[44][14] = 8'd14;
        rom[44][15] = 8'd5;
        rom[44][16] = -8'd65;
        rom[44][17] = 8'd11;
        rom[44][18] = -8'd51;
        rom[44][19] = -8'd26;
        rom[44][20] = 8'd4;
        rom[44][21] = -8'd6;
        rom[44][22] = -8'd14;
        rom[44][23] = -8'd7;
        rom[44][24] = -8'd13;
        rom[44][25] = 8'd17;
        rom[44][26] = 8'd35;
        rom[44][27] = 8'd15;
        rom[44][28] = -8'd27;
        rom[44][29] = 8'd19;
        rom[44][30] = 8'd3;
        rom[44][31] = -8'd9;
        rom[44][32] = -8'd3;
        rom[44][33] = -8'd63;
        rom[44][34] = -8'd23;
        rom[44][35] = -8'd19;
        rom[44][36] = 8'd30;
        rom[44][37] = 8'd1;
        rom[44][38] = -8'd29;
        rom[44][39] = -8'd7;
        rom[44][40] = -8'd95;
        rom[44][41] = -8'd2;
        rom[44][42] = -8'd19;
        rom[44][43] = -8'd24;
        rom[44][44] = 8'd7;
        rom[44][45] = 8'd11;
        rom[44][46] = -8'd20;
        rom[44][47] = -8'd45;
        rom[44][48] = 8'd2;
        rom[44][49] = -8'd42;
        rom[44][50] = 8'd9;
        rom[44][51] = 8'd15;
        rom[44][52] = -8'd10;
        rom[44][53] = -8'd47;
        rom[44][54] = -8'd22;
        rom[44][55] = 8'd12;
        rom[44][56] = 8'd35;
        rom[44][57] = 8'd2;
        rom[44][58] = 8'd3;
        rom[44][59] = -8'd34;
        rom[44][60] = 8'd11;
        rom[44][61] = -8'd3;
        rom[44][62] = -8'd41;
        rom[44][63] = -8'd19;
        rom[45][0] = 8'd13;
        rom[45][1] = -8'd9;
        rom[45][2] = 8'd8;
        rom[45][3] = -8'd12;
        rom[45][4] = 8'd8;
        rom[45][5] = 8'd16;
        rom[45][6] = -8'd9;
        rom[45][7] = -8'd8;
        rom[45][8] = -8'd16;
        rom[45][9] = 8'd15;
        rom[45][10] = -8'd15;
        rom[45][11] = 8'd0;
        rom[45][12] = 8'd36;
        rom[45][13] = -8'd58;
        rom[45][14] = -8'd5;
        rom[45][15] = 8'd0;
        rom[45][16] = 8'd25;
        rom[45][17] = 8'd11;
        rom[45][18] = -8'd23;
        rom[45][19] = 8'd60;
        rom[45][20] = 8'd4;
        rom[45][21] = 8'd68;
        rom[45][22] = 8'd46;
        rom[45][23] = -8'd4;
        rom[45][24] = 8'd20;
        rom[45][25] = 8'd9;
        rom[45][26] = -8'd34;
        rom[45][27] = 8'd13;
        rom[45][28] = 8'd4;
        rom[45][29] = -8'd14;
        rom[45][30] = 8'd42;
        rom[45][31] = -8'd2;
        rom[45][32] = 8'd14;
        rom[45][33] = -8'd15;
        rom[45][34] = 8'd17;
        rom[45][35] = 8'd0;
        rom[45][36] = 8'd30;
        rom[45][37] = 8'd23;
        rom[45][38] = 8'd20;
        rom[45][39] = -8'd27;
        rom[45][40] = -8'd17;
        rom[45][41] = 8'd19;
        rom[45][42] = 8'd24;
        rom[45][43] = -8'd15;
        rom[45][44] = 8'd2;
        rom[45][45] = 8'd15;
        rom[45][46] = 8'd38;
        rom[45][47] = 8'd12;
        rom[45][48] = 8'd23;
        rom[45][49] = 8'd0;
        rom[45][50] = 8'd18;
        rom[45][51] = -8'd14;
        rom[45][52] = 8'd30;
        rom[45][53] = 8'd6;
        rom[45][54] = 8'd7;
        rom[45][55] = -8'd18;
        rom[45][56] = -8'd13;
        rom[45][57] = -8'd29;
        rom[45][58] = 8'd10;
        rom[45][59] = 8'd56;
        rom[45][60] = 8'd26;
        rom[45][61] = 8'd17;
        rom[45][62] = 8'd12;
        rom[45][63] = 8'd41;
        rom[46][0] = 8'd1;
        rom[46][1] = -8'd13;
        rom[46][2] = 8'd15;
        rom[46][3] = 8'd3;
        rom[46][4] = 8'd2;
        rom[46][5] = 8'd17;
        rom[46][6] = -8'd31;
        rom[46][7] = 8'd3;
        rom[46][8] = -8'd82;
        rom[46][9] = -8'd25;
        rom[46][10] = -8'd49;
        rom[46][11] = -8'd29;
        rom[46][12] = -8'd21;
        rom[46][13] = 8'd31;
        rom[46][14] = -8'd4;
        rom[46][15] = -8'd49;
        rom[46][16] = -8'd14;
        rom[46][17] = 8'd37;
        rom[46][18] = -8'd26;
        rom[46][19] = 8'd2;
        rom[46][20] = -8'd11;
        rom[46][21] = -8'd5;
        rom[46][22] = -8'd25;
        rom[46][23] = 8'd24;
        rom[46][24] = -8'd3;
        rom[46][25] = -8'd84;
        rom[46][26] = 8'd34;
        rom[46][27] = 8'd24;
        rom[46][28] = -8'd40;
        rom[46][29] = -8'd43;
        rom[46][30] = 8'd13;
        rom[46][31] = 8'd5;
        rom[46][32] = 8'd5;
        rom[46][33] = -8'd9;
        rom[46][34] = -8'd8;
        rom[46][35] = -8'd12;
        rom[46][36] = 8'd2;
        rom[46][37] = 8'd2;
        rom[46][38] = 8'd2;
        rom[46][39] = -8'd19;
        rom[46][40] = 8'd3;
        rom[46][41] = 8'd42;
        rom[46][42] = -8'd14;
        rom[46][43] = 8'd35;
        rom[46][44] = -8'd37;
        rom[46][45] = 8'd34;
        rom[46][46] = -8'd15;
        rom[46][47] = -8'd9;
        rom[46][48] = -8'd1;
        rom[46][49] = 8'd17;
        rom[46][50] = -8'd7;
        rom[46][51] = 8'd26;
        rom[46][52] = 8'd22;
        rom[46][53] = -8'd23;
        rom[46][54] = -8'd32;
        rom[46][55] = -8'd52;
        rom[46][56] = 8'd6;
        rom[46][57] = 8'd0;
        rom[46][58] = -8'd1;
        rom[46][59] = 8'd6;
        rom[46][60] = -8'd54;
        rom[46][61] = -8'd16;
        rom[46][62] = 8'd34;
        rom[46][63] = -8'd31;
        rom[47][0] = 8'd12;
        rom[47][1] = 8'd38;
        rom[47][2] = -8'd32;
        rom[47][3] = -8'd3;
        rom[47][4] = 8'd34;
        rom[47][5] = -8'd24;
        rom[47][6] = 8'd4;
        rom[47][7] = 8'd17;
        rom[47][8] = 8'd27;
        rom[47][9] = -8'd21;
        rom[47][10] = 8'd21;
        rom[47][11] = 8'd57;
        rom[47][12] = -8'd32;
        rom[47][13] = -8'd8;
        rom[47][14] = 8'd28;
        rom[47][15] = -8'd2;
        rom[47][16] = 8'd57;
        rom[47][17] = 8'd42;
        rom[47][18] = -8'd7;
        rom[47][19] = -8'd14;
        rom[47][20] = 8'd7;
        rom[47][21] = 8'd28;
        rom[47][22] = 8'd21;
        rom[47][23] = -8'd37;
        rom[47][24] = -8'd37;
        rom[47][25] = -8'd3;
        rom[47][26] = 8'd1;
        rom[47][27] = 8'd41;
        rom[47][28] = -8'd40;
        rom[47][29] = 8'd22;
        rom[47][30] = -8'd31;
        rom[47][31] = 8'd14;
        rom[47][32] = -8'd38;
        rom[47][33] = 8'd38;
        rom[47][34] = -8'd10;
        rom[47][35] = 8'd52;
        rom[47][36] = -8'd37;
        rom[47][37] = 8'd16;
        rom[47][38] = 8'd9;
        rom[47][39] = 8'd14;
        rom[47][40] = -8'd1;
        rom[47][41] = -8'd26;
        rom[47][42] = 8'd17;
        rom[47][43] = -8'd21;
        rom[47][44] = 8'd52;
        rom[47][45] = 8'd54;
        rom[47][46] = 8'd28;
        rom[47][47] = 8'd2;
        rom[47][48] = 8'd50;
        rom[47][49] = 8'd44;
        rom[47][50] = -8'd14;
        rom[47][51] = 8'd60;
        rom[47][52] = -8'd32;
        rom[47][53] = 8'd46;
        rom[47][54] = -8'd30;
        rom[47][55] = -8'd30;
        rom[47][56] = -8'd25;
        rom[47][57] = 8'd19;
        rom[47][58] = 8'd5;
        rom[47][59] = 8'd70;
        rom[47][60] = -8'd24;
        rom[47][61] = -8'd19;
        rom[47][62] = -8'd19;
        rom[47][63] = -8'd45;
        rom[48][0] = -8'd12;
        rom[48][1] = 8'd23;
        rom[48][2] = -8'd34;
        rom[48][3] = 8'd16;
        rom[48][4] = 8'd3;
        rom[48][5] = -8'd10;
        rom[48][6] = -8'd41;
        rom[48][7] = -8'd36;
        rom[48][8] = 8'd15;
        rom[48][9] = -8'd13;
        rom[48][10] = -8'd7;
        rom[48][11] = 8'd7;
        rom[48][12] = -8'd13;
        rom[48][13] = -8'd5;
        rom[48][14] = -8'd5;
        rom[48][15] = -8'd12;
        rom[48][16] = 8'd25;
        rom[48][17] = -8'd32;
        rom[48][18] = -8'd54;
        rom[48][19] = 8'd24;
        rom[48][20] = -8'd2;
        rom[48][21] = 8'd28;
        rom[48][22] = -8'd15;
        rom[48][23] = 8'd7;
        rom[48][24] = -8'd52;
        rom[48][25] = 8'd16;
        rom[48][26] = -8'd46;
        rom[48][27] = -8'd9;
        rom[48][28] = -8'd4;
        rom[48][29] = -8'd8;
        rom[48][30] = 8'd0;
        rom[48][31] = 8'd22;
        rom[48][32] = -8'd33;
        rom[48][33] = -8'd20;
        rom[48][34] = 8'd10;
        rom[48][35] = -8'd1;
        rom[48][36] = -8'd23;
        rom[48][37] = 8'd3;
        rom[48][38] = 8'd26;
        rom[48][39] = 8'd11;
        rom[48][40] = 8'd12;
        rom[48][41] = 8'd8;
        rom[48][42] = -8'd46;
        rom[48][43] = 8'd21;
        rom[48][44] = -8'd33;
        rom[48][45] = 8'd7;
        rom[48][46] = 8'd0;
        rom[48][47] = 8'd4;
        rom[48][48] = -8'd50;
        rom[48][49] = -8'd24;
        rom[48][50] = 8'd25;
        rom[48][51] = 8'd12;
        rom[48][52] = -8'd45;
        rom[48][53] = -8'd40;
        rom[48][54] = -8'd52;
        rom[48][55] = 8'd21;
        rom[48][56] = 8'd28;
        rom[48][57] = -8'd61;
        rom[48][58] = -8'd10;
        rom[48][59] = 8'd42;
        rom[48][60] = -8'd39;
        rom[48][61] = 8'd9;
        rom[48][62] = -8'd36;
        rom[48][63] = 8'd14;
        rom[49][0] = -8'd22;
        rom[49][1] = 8'd17;
        rom[49][2] = 8'd37;
        rom[49][3] = -8'd33;
        rom[49][4] = -8'd13;
        rom[49][5] = 8'd12;
        rom[49][6] = -8'd51;
        rom[49][7] = -8'd25;
        rom[49][8] = 8'd17;
        rom[49][9] = 8'd29;
        rom[49][10] = 8'd31;
        rom[49][11] = 8'd13;
        rom[49][12] = 8'd68;
        rom[49][13] = 8'd1;
        rom[49][14] = 8'd1;
        rom[49][15] = -8'd12;
        rom[49][16] = 8'd13;
        rom[49][17] = -8'd25;
        rom[49][18] = -8'd24;
        rom[49][19] = 8'd64;
        rom[49][20] = -8'd10;
        rom[49][21] = -8'd53;
        rom[49][22] = 8'd65;
        rom[49][23] = -8'd32;
        rom[49][24] = -8'd25;
        rom[49][25] = -8'd27;
        rom[49][26] = -8'd11;
        rom[49][27] = -8'd11;
        rom[49][28] = 8'd21;
        rom[49][29] = -8'd16;
        rom[49][30] = 8'd49;
        rom[49][31] = 8'd2;
        rom[49][32] = -8'd14;
        rom[49][33] = 8'd44;
        rom[49][34] = 8'd2;
        rom[49][35] = -8'd42;
        rom[49][36] = -8'd63;
        rom[49][37] = 8'd0;
        rom[49][38] = 8'd29;
        rom[49][39] = 8'd22;
        rom[49][40] = -8'd18;
        rom[49][41] = -8'd7;
        rom[49][42] = 8'd47;
        rom[49][43] = -8'd4;
        rom[49][44] = -8'd40;
        rom[49][45] = 8'd1;
        rom[49][46] = -8'd10;
        rom[49][47] = 8'd6;
        rom[49][48] = -8'd13;
        rom[49][49] = 8'd14;
        rom[49][50] = -8'd17;
        rom[49][51] = -8'd18;
        rom[49][52] = 8'd3;
        rom[49][53] = 8'd39;
        rom[49][54] = 8'd19;
        rom[49][55] = -8'd19;
        rom[49][56] = 8'd1;
        rom[49][57] = -8'd17;
        rom[49][58] = 8'd3;
        rom[49][59] = -8'd9;
        rom[49][60] = 8'd3;
        rom[49][61] = -8'd13;
        rom[49][62] = -8'd29;
        rom[49][63] = 8'd17;
        rom[50][0] = 8'd17;
        rom[50][1] = -8'd27;
        rom[50][2] = 8'd1;
        rom[50][3] = -8'd2;
        rom[50][4] = -8'd26;
        rom[50][5] = 8'd2;
        rom[50][6] = 8'd16;
        rom[50][7] = -8'd29;
        rom[50][8] = -8'd29;
        rom[50][9] = 8'd9;
        rom[50][10] = -8'd28;
        rom[50][11] = -8'd43;
        rom[50][12] = 8'd18;
        rom[50][13] = -8'd24;
        rom[50][14] = -8'd21;
        rom[50][15] = -8'd34;
        rom[50][16] = -8'd24;
        rom[50][17] = 8'd5;
        rom[50][18] = 8'd5;
        rom[50][19] = -8'd36;
        rom[50][20] = -8'd12;
        rom[50][21] = -8'd3;
        rom[50][22] = -8'd46;
        rom[50][23] = -8'd36;
        rom[50][24] = 8'd10;
        rom[50][25] = -8'd13;
        rom[50][26] = 8'd27;
        rom[50][27] = -8'd49;
        rom[50][28] = -8'd2;
        rom[50][29] = 8'd0;
        rom[50][30] = 8'd0;
        rom[50][31] = -8'd68;
        rom[50][32] = -8'd10;
        rom[50][33] = 8'd11;
        rom[50][34] = -8'd15;
        rom[50][35] = -8'd12;
        rom[50][36] = 8'd25;
        rom[50][37] = -8'd13;
        rom[50][38] = -8'd8;
        rom[50][39] = -8'd36;
        rom[50][40] = -8'd14;
        rom[50][41] = -8'd24;
        rom[50][42] = -8'd15;
        rom[50][43] = -8'd6;
        rom[50][44] = -8'd14;
        rom[50][45] = -8'd6;
        rom[50][46] = 8'd4;
        rom[50][47] = -8'd37;
        rom[50][48] = -8'd27;
        rom[50][49] = 8'd6;
        rom[50][50] = -8'd12;
        rom[50][51] = -8'd66;
        rom[50][52] = 8'd19;
        rom[50][53] = 8'd0;
        rom[50][54] = 8'd20;
        rom[50][55] = -8'd27;
        rom[50][56] = -8'd3;
        rom[50][57] = -8'd38;
        rom[50][58] = 8'd26;
        rom[50][59] = -8'd13;
        rom[50][60] = -8'd2;
        rom[50][61] = 8'd14;
        rom[50][62] = 8'd58;
        rom[50][63] = -8'd30;
        rom[51][0] = 8'd33;
        rom[51][1] = -8'd4;
        rom[51][2] = 8'd34;
        rom[51][3] = 8'd12;
        rom[51][4] = 8'd8;
        rom[51][5] = 8'd12;
        rom[51][6] = 8'd34;
        rom[51][7] = 8'd25;
        rom[51][8] = -8'd4;
        rom[51][9] = -8'd13;
        rom[51][10] = 8'd0;
        rom[51][11] = -8'd30;
        rom[51][12] = 8'd44;
        rom[51][13] = -8'd38;
        rom[51][14] = -8'd54;
        rom[51][15] = 8'd19;
        rom[51][16] = 8'd12;
        rom[51][17] = -8'd12;
        rom[51][18] = -8'd17;
        rom[51][19] = 8'd35;
        rom[51][20] = -8'd5;
        rom[51][21] = -8'd13;
        rom[51][22] = -8'd49;
        rom[51][23] = -8'd10;
        rom[51][24] = 8'd12;
        rom[51][25] = 8'd9;
        rom[51][26] = -8'd17;
        rom[51][27] = -8'd30;
        rom[51][28] = -8'd21;
        rom[51][29] = -8'd42;
        rom[51][30] = -8'd20;
        rom[51][31] = -8'd18;
        rom[51][32] = 8'd5;
        rom[51][33] = 8'd39;
        rom[51][34] = -8'd68;
        rom[51][35] = -8'd8;
        rom[51][36] = 8'd34;
        rom[51][37] = 8'd20;
        rom[51][38] = 8'd25;
        rom[51][39] = -8'd6;
        rom[51][40] = -8'd9;
        rom[51][41] = 8'd5;
        rom[51][42] = 8'd7;
        rom[51][43] = -8'd48;
        rom[51][44] = 8'd2;
        rom[51][45] = -8'd3;
        rom[51][46] = 8'd8;
        rom[51][47] = 8'd19;
        rom[51][48] = 8'd23;
        rom[51][49] = -8'd14;
        rom[51][50] = -8'd28;
        rom[51][51] = -8'd27;
        rom[51][52] = -8'd8;
        rom[51][53] = -8'd35;
        rom[51][54] = -8'd36;
        rom[51][55] = -8'd6;
        rom[51][56] = -8'd15;
        rom[51][57] = 8'd11;
        rom[51][58] = 8'd4;
        rom[51][59] = 8'd4;
        rom[51][60] = 8'd26;
        rom[51][61] = -8'd4;
        rom[51][62] = 8'd13;
        rom[51][63] = 8'd10;
        rom[52][0] = 8'd3;
        rom[52][1] = -8'd26;
        rom[52][2] = 8'd35;
        rom[52][3] = 8'd1;
        rom[52][4] = 8'd26;
        rom[52][5] = -8'd16;
        rom[52][6] = -8'd8;
        rom[52][7] = -8'd8;
        rom[52][8] = 8'd18;
        rom[52][9] = -8'd13;
        rom[52][10] = 8'd0;
        rom[52][11] = 8'd3;
        rom[52][12] = -8'd39;
        rom[52][13] = -8'd2;
        rom[52][14] = 8'd51;
        rom[52][15] = 8'd54;
        rom[52][16] = -8'd35;
        rom[52][17] = 8'd23;
        rom[52][18] = 8'd15;
        rom[52][19] = -8'd18;
        rom[52][20] = 8'd4;
        rom[52][21] = 8'd18;
        rom[52][22] = 8'd46;
        rom[52][23] = -8'd24;
        rom[52][24] = -8'd16;
        rom[52][25] = 8'd4;
        rom[52][26] = 8'd10;
        rom[52][27] = 8'd11;
        rom[52][28] = -8'd4;
        rom[52][29] = 8'd9;
        rom[52][30] = 8'd0;
        rom[52][31] = -8'd3;
        rom[52][32] = -8'd45;
        rom[52][33] = -8'd37;
        rom[52][34] = -8'd2;
        rom[52][35] = 8'd11;
        rom[52][36] = -8'd83;
        rom[52][37] = -8'd39;
        rom[52][38] = -8'd24;
        rom[52][39] = -8'd6;
        rom[52][40] = 8'd27;
        rom[52][41] = 8'd29;
        rom[52][42] = -8'd20;
        rom[52][43] = -8'd8;
        rom[52][44] = -8'd30;
        rom[52][45] = -8'd9;
        rom[52][46] = -8'd22;
        rom[52][47] = 8'd3;
        rom[52][48] = 8'd27;
        rom[52][49] = -8'd3;
        rom[52][50] = 8'd9;
        rom[52][51] = 8'd6;
        rom[52][52] = 8'd59;
        rom[52][53] = 8'd6;
        rom[52][54] = 8'd3;
        rom[52][55] = 8'd13;
        rom[52][56] = -8'd27;
        rom[52][57] = 8'd8;
        rom[52][58] = 8'd15;
        rom[52][59] = 8'd15;
        rom[52][60] = -8'd13;
        rom[52][61] = -8'd7;
        rom[52][62] = -8'd27;
        rom[52][63] = 8'd19;
        rom[53][0] = -8'd5;
        rom[53][1] = 8'd23;
        rom[53][2] = -8'd10;
        rom[53][3] = 8'd2;
        rom[53][4] = -8'd28;
        rom[53][5] = 8'd7;
        rom[53][6] = -8'd52;
        rom[53][7] = 8'd9;
        rom[53][8] = -8'd25;
        rom[53][9] = -8'd1;
        rom[53][10] = -8'd32;
        rom[53][11] = 8'd19;
        rom[53][12] = 8'd14;
        rom[53][13] = 8'd4;
        rom[53][14] = 8'd19;
        rom[53][15] = 8'd17;
        rom[53][16] = 8'd42;
        rom[53][17] = 8'd7;
        rom[53][18] = 8'd20;
        rom[53][19] = 8'd25;
        rom[53][20] = -8'd4;
        rom[53][21] = -8'd3;
        rom[53][22] = 8'd2;
        rom[53][23] = -8'd6;
        rom[53][24] = 8'd0;
        rom[53][25] = -8'd45;
        rom[53][26] = -8'd5;
        rom[53][27] = 8'd22;
        rom[53][28] = 8'd7;
        rom[53][29] = -8'd31;
        rom[53][30] = 8'd2;
        rom[53][31] = -8'd11;
        rom[53][32] = -8'd41;
        rom[53][33] = -8'd36;
        rom[53][34] = 8'd14;
        rom[53][35] = -8'd19;
        rom[53][36] = 8'd6;
        rom[53][37] = 8'd9;
        rom[53][38] = 8'd36;
        rom[53][39] = 8'd0;
        rom[53][40] = -8'd31;
        rom[53][41] = -8'd30;
        rom[53][42] = -8'd21;
        rom[53][43] = -8'd26;
        rom[53][44] = -8'd20;
        rom[53][45] = 8'd27;
        rom[53][46] = -8'd31;
        rom[53][47] = 8'd34;
        rom[53][48] = -8'd5;
        rom[53][49] = -8'd40;
        rom[53][50] = 8'd33;
        rom[53][51] = -8'd26;
        rom[53][52] = -8'd23;
        rom[53][53] = -8'd36;
        rom[53][54] = 8'd35;
        rom[53][55] = -8'd25;
        rom[53][56] = 8'd12;
        rom[53][57] = 8'd8;
        rom[53][58] = -8'd8;
        rom[53][59] = 8'd26;
        rom[53][60] = 8'd10;
        rom[53][61] = -8'd15;
        rom[53][62] = 8'd10;
        rom[53][63] = -8'd35;
        rom[54][0] = -8'd2;
        rom[54][1] = 8'd3;
        rom[54][2] = 8'd5;
        rom[54][3] = -8'd2;
        rom[54][4] = 8'd8;
        rom[54][5] = 8'd8;
        rom[54][6] = -8'd4;
        rom[54][7] = 8'd0;
        rom[54][8] = 8'd3;
        rom[54][9] = -8'd9;
        rom[54][10] = -8'd5;
        rom[54][11] = 8'd1;
        rom[54][12] = 8'd0;
        rom[54][13] = 8'd2;
        rom[54][14] = 8'd4;
        rom[54][15] = -8'd6;
        rom[54][16] = -8'd1;
        rom[54][17] = 8'd12;
        rom[54][18] = 8'd7;
        rom[54][19] = 8'd5;
        rom[54][20] = 8'd5;
        rom[54][21] = -8'd6;
        rom[54][22] = 8'd5;
        rom[54][23] = 8'd9;
        rom[54][24] = -8'd3;
        rom[54][25] = 8'd3;
        rom[54][26] = 8'd4;
        rom[54][27] = -8'd1;
        rom[54][28] = 8'd6;
        rom[54][29] = -8'd2;
        rom[54][30] = -8'd4;
        rom[54][31] = 8'd10;
        rom[54][32] = 8'd7;
        rom[54][33] = -8'd5;
        rom[54][34] = 8'd4;
        rom[54][35] = 8'd0;
        rom[54][36] = 8'd7;
        rom[54][37] = -8'd7;
        rom[54][38] = -8'd2;
        rom[54][39] = -8'd11;
        rom[54][40] = 8'd9;
        rom[54][41] = 8'd0;
        rom[54][42] = -8'd7;
        rom[54][43] = 8'd3;
        rom[54][44] = 8'd6;
        rom[54][45] = -8'd13;
        rom[54][46] = -8'd7;
        rom[54][47] = 8'd11;
        rom[54][48] = 8'd6;
        rom[54][49] = -8'd7;
        rom[54][50] = 8'd4;
        rom[54][51] = -8'd6;
        rom[54][52] = 8'd6;
        rom[54][53] = -8'd2;
        rom[54][54] = 8'd11;
        rom[54][55] = -8'd12;
        rom[54][56] = -8'd1;
        rom[54][57] = 8'd1;
        rom[54][58] = 8'd4;
        rom[54][59] = 8'd10;
        rom[54][60] = 8'd2;
        rom[54][61] = -8'd3;
        rom[54][62] = 8'd7;
        rom[54][63] = -8'd5;
        rom[55][0] = -8'd22;
        rom[55][1] = -8'd13;
        rom[55][2] = -8'd13;
        rom[55][3] = 8'd15;
        rom[55][4] = -8'd20;
        rom[55][5] = 8'd0;
        rom[55][6] = -8'd29;
        rom[55][7] = 8'd19;
        rom[55][8] = 8'd37;
        rom[55][9] = 8'd5;
        rom[55][10] = 8'd6;
        rom[55][11] = -8'd42;
        rom[55][12] = -8'd36;
        rom[55][13] = 8'd43;
        rom[55][14] = -8'd46;
        rom[55][15] = 8'd40;
        rom[55][16] = -8'd30;
        rom[55][17] = 8'd32;
        rom[55][18] = -8'd13;
        rom[55][19] = 8'd14;
        rom[55][20] = -8'd6;
        rom[55][21] = 8'd3;
        rom[55][22] = -8'd20;
        rom[55][23] = 8'd6;
        rom[55][24] = -8'd56;
        rom[55][25] = -8'd1;
        rom[55][26] = -8'd12;
        rom[55][27] = -8'd60;
        rom[55][28] = -8'd3;
        rom[55][29] = -8'd13;
        rom[55][30] = 8'd67;
        rom[55][31] = 8'd34;
        rom[55][32] = -8'd27;
        rom[55][33] = 8'd7;
        rom[55][34] = 8'd3;
        rom[55][35] = 8'd4;
        rom[55][36] = -8'd16;
        rom[55][37] = 8'd1;
        rom[55][38] = -8'd17;
        rom[55][39] = 8'd13;
        rom[55][40] = 8'd49;
        rom[55][41] = 8'd38;
        rom[55][42] = 8'd2;
        rom[55][43] = 8'd0;
        rom[55][44] = -8'd7;
        rom[55][45] = -8'd47;
        rom[55][46] = -8'd30;
        rom[55][47] = -8'd31;
        rom[55][48] = -8'd2;
        rom[55][49] = 8'd26;
        rom[55][50] = -8'd41;
        rom[55][51] = 8'd15;
        rom[55][52] = 8'd28;
        rom[55][53] = -8'd1;
        rom[55][54] = 8'd1;
        rom[55][55] = 8'd30;
        rom[55][56] = 8'd9;
        rom[55][57] = 8'd31;
        rom[55][58] = -8'd6;
        rom[55][59] = -8'd9;
        rom[55][60] = -8'd11;
        rom[55][61] = 8'd5;
        rom[55][62] = 8'd10;
        rom[55][63] = 8'd3;
        rom[56][0] = -8'd37;
        rom[56][1] = 8'd14;
        rom[56][2] = 8'd23;
        rom[56][3] = -8'd49;
        rom[56][4] = -8'd27;
        rom[56][5] = -8'd19;
        rom[56][6] = -8'd8;
        rom[56][7] = -8'd11;
        rom[56][8] = 8'd6;
        rom[56][9] = -8'd7;
        rom[56][10] = -8'd5;
        rom[56][11] = -8'd58;
        rom[56][12] = -8'd56;
        rom[56][13] = 8'd2;
        rom[56][14] = 8'd11;
        rom[56][15] = -8'd24;
        rom[56][16] = 8'd40;
        rom[56][17] = -8'd1;
        rom[56][18] = 8'd3;
        rom[56][19] = 8'd13;
        rom[56][20] = -8'd8;
        rom[56][21] = 8'd1;
        rom[56][22] = 8'd23;
        rom[56][23] = -8'd25;
        rom[56][24] = -8'd82;
        rom[56][25] = -8'd8;
        rom[56][26] = 8'd47;
        rom[56][27] = 8'd28;
        rom[56][28] = 8'd7;
        rom[56][29] = 8'd19;
        rom[56][30] = 8'd11;
        rom[56][31] = 8'd9;
        rom[56][32] = -8'd37;
        rom[56][33] = -8'd48;
        rom[56][34] = -8'd15;
        rom[56][35] = -8'd3;
        rom[56][36] = -8'd29;
        rom[56][37] = -8'd6;
        rom[56][38] = -8'd18;
        rom[56][39] = 8'd27;
        rom[56][40] = 8'd14;
        rom[56][41] = -8'd32;
        rom[56][42] = -8'd40;
        rom[56][43] = -8'd2;
        rom[56][44] = -8'd15;
        rom[56][45] = -8'd32;
        rom[56][46] = 8'd0;
        rom[56][47] = -8'd46;
        rom[56][48] = -8'd45;
        rom[56][49] = 8'd12;
        rom[56][50] = 8'd28;
        rom[56][51] = 8'd14;
        rom[56][52] = 8'd1;
        rom[56][53] = 8'd7;
        rom[56][54] = -8'd1;
        rom[56][55] = -8'd14;
        rom[56][56] = 8'd16;
        rom[56][57] = -8'd1;
        rom[56][58] = -8'd19;
        rom[56][59] = -8'd40;
        rom[56][60] = -8'd3;
        rom[56][61] = 8'd31;
        rom[56][62] = -8'd17;
        rom[56][63] = -8'd26;
        rom[57][0] = 8'd24;
        rom[57][1] = -8'd21;
        rom[57][2] = -8'd13;
        rom[57][3] = 8'd23;
        rom[57][4] = -8'd2;
        rom[57][5] = 8'd26;
        rom[57][6] = 8'd16;
        rom[57][7] = 8'd18;
        rom[57][8] = 8'd15;
        rom[57][9] = -8'd10;
        rom[57][10] = 8'd26;
        rom[57][11] = -8'd69;
        rom[57][12] = -8'd31;
        rom[57][13] = -8'd16;
        rom[57][14] = -8'd42;
        rom[57][15] = -8'd8;
        rom[57][16] = -8'd10;
        rom[57][17] = 8'd18;
        rom[57][18] = -8'd63;
        rom[57][19] = 8'd69;
        rom[57][20] = 8'd0;
        rom[57][21] = 8'd30;
        rom[57][22] = -8'd7;
        rom[57][23] = 8'd22;
        rom[57][24] = 8'd34;
        rom[57][25] = -8'd14;
        rom[57][26] = 8'd0;
        rom[57][27] = -8'd23;
        rom[57][28] = 8'd2;
        rom[57][29] = 8'd36;
        rom[57][30] = -8'd44;
        rom[57][31] = 8'd5;
        rom[57][32] = 8'd60;
        rom[57][33] = -8'd11;
        rom[57][34] = -8'd8;
        rom[57][35] = -8'd23;
        rom[57][36] = 8'd0;
        rom[57][37] = 8'd38;
        rom[57][38] = 8'd66;
        rom[57][39] = -8'd7;
        rom[57][40] = -8'd39;
        rom[57][41] = -8'd5;
        rom[57][42] = 8'd13;
        rom[57][43] = 8'd22;
        rom[57][44] = 8'd4;
        rom[57][45] = -8'd20;
        rom[57][46] = -8'd14;
        rom[57][47] = 8'd32;
        rom[57][48] = 8'd11;
        rom[57][49] = -8'd12;
        rom[57][50] = -8'd38;
        rom[57][51] = -8'd12;
        rom[57][52] = 8'd3;
        rom[57][53] = -8'd54;
        rom[57][54] = 8'd18;
        rom[57][55] = 8'd8;
        rom[57][56] = 8'd25;
        rom[57][57] = 8'd26;
        rom[57][58] = -8'd5;
        rom[57][59] = 8'd20;
        rom[57][60] = 8'd29;
        rom[57][61] = -8'd34;
        rom[57][62] = -8'd5;
        rom[57][63] = -8'd33;
        rom[58][0] = -8'd1;
        rom[58][1] = 8'd14;
        rom[58][2] = -8'd15;
        rom[58][3] = 8'd12;
        rom[58][4] = 8'd7;
        rom[58][5] = 8'd30;
        rom[58][6] = -8'd20;
        rom[58][7] = 8'd43;
        rom[58][8] = -8'd20;
        rom[58][9] = 8'd12;
        rom[58][10] = 8'd46;
        rom[58][11] = -8'd38;
        rom[58][12] = -8'd28;
        rom[58][13] = -8'd27;
        rom[58][14] = -8'd12;
        rom[58][15] = 8'd40;
        rom[58][16] = 8'd68;
        rom[58][17] = 8'd50;
        rom[58][18] = -8'd85;
        rom[58][19] = 8'd6;
        rom[58][20] = 8'd0;
        rom[58][21] = -8'd30;
        rom[58][22] = 8'd11;
        rom[58][23] = -8'd15;
        rom[58][24] = 8'd30;
        rom[58][25] = 8'd14;
        rom[58][26] = 8'd49;
        rom[58][27] = 8'd28;
        rom[58][28] = -8'd4;
        rom[58][29] = -8'd39;
        rom[58][30] = -8'd35;
        rom[58][31] = 8'd15;
        rom[58][32] = -8'd7;
        rom[58][33] = -8'd14;
        rom[58][34] = -8'd24;
        rom[58][35] = -8'd73;
        rom[58][36] = -8'd22;
        rom[58][37] = 8'd18;
        rom[58][38] = 8'd23;
        rom[58][39] = -8'd26;
        rom[58][40] = 8'd3;
        rom[58][41] = -8'd2;
        rom[58][42] = -8'd13;
        rom[58][43] = -8'd2;
        rom[58][44] = -8'd25;
        rom[58][45] = -8'd19;
        rom[58][46] = 8'd11;
        rom[58][47] = -8'd18;
        rom[58][48] = -8'd23;
        rom[58][49] = -8'd58;
        rom[58][50] = -8'd15;
        rom[58][51] = -8'd106;
        rom[58][52] = 8'd2;
        rom[58][53] = -8'd16;
        rom[58][54] = -8'd51;
        rom[58][55] = -8'd5;
        rom[58][56] = 8'd2;
        rom[58][57] = 8'd12;
        rom[58][58] = 8'd23;
        rom[58][59] = -8'd3;
        rom[58][60] = 8'd64;
        rom[58][61] = 8'd39;
        rom[58][62] = -8'd30;
        rom[58][63] = 8'd0;
        rom[59][0] = 8'd21;
        rom[59][1] = 8'd11;
        rom[59][2] = -8'd19;
        rom[59][3] = -8'd23;
        rom[59][4] = -8'd13;
        rom[59][5] = -8'd14;
        rom[59][6] = -8'd2;
        rom[59][7] = 8'd31;
        rom[59][8] = 8'd24;
        rom[59][9] = 8'd18;
        rom[59][10] = 8'd17;
        rom[59][11] = -8'd3;
        rom[59][12] = -8'd27;
        rom[59][13] = -8'd10;
        rom[59][14] = 8'd3;
        rom[59][15] = 8'd15;
        rom[59][16] = -8'd42;
        rom[59][17] = 8'd33;
        rom[59][18] = 8'd40;
        rom[59][19] = 8'd14;
        rom[59][20] = -8'd7;
        rom[59][21] = 8'd1;
        rom[59][22] = 8'd23;
        rom[59][23] = 8'd5;
        rom[59][24] = -8'd31;
        rom[59][25] = -8'd22;
        rom[59][26] = -8'd11;
        rom[59][27] = 8'd3;
        rom[59][28] = -8'd25;
        rom[59][29] = 8'd13;
        rom[59][30] = -8'd27;
        rom[59][31] = 8'd14;
        rom[59][32] = -8'd52;
        rom[59][33] = 8'd10;
        rom[59][34] = 8'd33;
        rom[59][35] = 8'd18;
        rom[59][36] = 8'd9;
        rom[59][37] = -8'd12;
        rom[59][38] = -8'd13;
        rom[59][39] = -8'd13;
        rom[59][40] = -8'd5;
        rom[59][41] = -8'd9;
        rom[59][42] = -8'd3;
        rom[59][43] = 8'd35;
        rom[59][44] = -8'd5;
        rom[59][45] = 8'd6;
        rom[59][46] = -8'd55;
        rom[59][47] = -8'd51;
        rom[59][48] = -8'd19;
        rom[59][49] = 8'd11;
        rom[59][50] = -8'd3;
        rom[59][51] = -8'd14;
        rom[59][52] = 8'd20;
        rom[59][53] = 8'd24;
        rom[59][54] = -8'd11;
        rom[59][55] = 8'd6;
        rom[59][56] = -8'd13;
        rom[59][57] = -8'd34;
        rom[59][58] = 8'd11;
        rom[59][59] = -8'd4;
        rom[59][60] = 8'd20;
        rom[59][61] = -8'd5;
        rom[59][62] = -8'd31;
        rom[59][63] = 8'd11;
        rom[60][0] = 8'd6;
        rom[60][1] = 8'd14;
        rom[60][2] = 8'd4;
        rom[60][3] = 8'd17;
        rom[60][4] = -8'd3;
        rom[60][5] = -8'd43;
        rom[60][6] = -8'd14;
        rom[60][7] = 8'd6;
        rom[60][8] = -8'd1;
        rom[60][9] = 8'd3;
        rom[60][10] = -8'd53;
        rom[60][11] = -8'd16;
        rom[60][12] = -8'd3;
        rom[60][13] = -8'd29;
        rom[60][14] = -8'd12;
        rom[60][15] = 8'd13;
        rom[60][16] = -8'd3;
        rom[60][17] = 8'd11;
        rom[60][18] = -8'd23;
        rom[60][19] = 8'd33;
        rom[60][20] = -8'd21;
        rom[60][21] = 8'd25;
        rom[60][22] = -8'd29;
        rom[60][23] = 8'd12;
        rom[60][24] = -8'd31;
        rom[60][25] = 8'd0;
        rom[60][26] = -8'd3;
        rom[60][27] = 8'd35;
        rom[60][28] = 8'd3;
        rom[60][29] = -8'd27;
        rom[60][30] = 8'd14;
        rom[60][31] = 8'd19;
        rom[60][32] = 8'd13;
        rom[60][33] = 8'd10;
        rom[60][34] = -8'd3;
        rom[60][35] = 8'd0;
        rom[60][36] = 8'd20;
        rom[60][37] = -8'd6;
        rom[60][38] = 8'd3;
        rom[60][39] = -8'd40;
        rom[60][40] = 8'd13;
        rom[60][41] = -8'd3;
        rom[60][42] = 8'd3;
        rom[60][43] = 8'd21;
        rom[60][44] = 8'd24;
        rom[60][45] = 8'd23;
        rom[60][46] = 8'd4;
        rom[60][47] = -8'd30;
        rom[60][48] = -8'd33;
        rom[60][49] = 8'd10;
        rom[60][50] = 8'd0;
        rom[60][51] = -8'd31;
        rom[60][52] = -8'd56;
        rom[60][53] = 8'd14;
        rom[60][54] = 8'd40;
        rom[60][55] = 8'd6;
        rom[60][56] = 8'd3;
        rom[60][57] = 8'd4;
        rom[60][58] = 8'd15;
        rom[60][59] = 8'd18;
        rom[60][60] = -8'd43;
        rom[60][61] = -8'd20;
        rom[60][62] = -8'd28;
        rom[60][63] = -8'd21;
        rom[61][0] = 8'd30;
        rom[61][1] = -8'd22;
        rom[61][2] = 8'd48;
        rom[61][3] = 8'd3;
        rom[61][4] = 8'd15;
        rom[61][5] = 8'd30;
        rom[61][6] = 8'd3;
        rom[61][7] = -8'd46;
        rom[61][8] = 8'd5;
        rom[61][9] = 8'd0;
        rom[61][10] = 8'd26;
        rom[61][11] = -8'd10;
        rom[61][12] = -8'd17;
        rom[61][13] = 8'd5;
        rom[61][14] = 8'd5;
        rom[61][15] = -8'd21;
        rom[61][16] = 8'd11;
        rom[61][17] = 8'd17;
        rom[61][18] = -8'd6;
        rom[61][19] = -8'd19;
        rom[61][20] = 8'd13;
        rom[61][21] = -8'd3;
        rom[61][22] = 8'd11;
        rom[61][23] = -8'd48;
        rom[61][24] = -8'd27;
        rom[61][25] = -8'd23;
        rom[61][26] = 8'd26;
        rom[61][27] = -8'd75;
        rom[61][28] = -8'd11;
        rom[61][29] = 8'd2;
        rom[61][30] = 8'd21;
        rom[61][31] = 8'd2;
        rom[61][32] = 8'd1;
        rom[61][33] = -8'd9;
        rom[61][34] = 8'd3;
        rom[61][35] = 8'd28;
        rom[61][36] = -8'd42;
        rom[61][37] = 8'd23;
        rom[61][38] = 8'd3;
        rom[61][39] = 8'd23;
        rom[61][40] = -8'd13;
        rom[61][41] = -8'd4;
        rom[61][42] = -8'd23;
        rom[61][43] = -8'd48;
        rom[61][44] = -8'd39;
        rom[61][45] = -8'd4;
        rom[61][46] = -8'd12;
        rom[61][47] = 8'd58;
        rom[61][48] = 8'd5;
        rom[61][49] = -8'd95;
        rom[61][50] = -8'd24;
        rom[61][51] = -8'd25;
        rom[61][52] = 8'd29;
        rom[61][53] = 8'd3;
        rom[61][54] = -8'd13;
        rom[61][55] = -8'd15;
        rom[61][56] = 8'd16;
        rom[61][57] = -8'd2;
        rom[61][58] = -8'd5;
        rom[61][59] = -8'd22;
        rom[61][60] = -8'd5;
        rom[61][61] = -8'd42;
        rom[61][62] = -8'd37;
        rom[61][63] = -8'd33;
        rom[62][0] = 8'd57;
        rom[62][1] = -8'd44;
        rom[62][2] = 8'd10;
        rom[62][3] = -8'd29;
        rom[62][4] = -8'd68;
        rom[62][5] = -8'd4;
        rom[62][6] = -8'd41;
        rom[62][7] = 8'd8;
        rom[62][8] = -8'd46;
        rom[62][9] = 8'd1;
        rom[62][10] = -8'd4;
        rom[62][11] = 8'd49;
        rom[62][12] = 8'd47;
        rom[62][13] = -8'd44;
        rom[62][14] = -8'd18;
        rom[62][15] = -8'd5;
        rom[62][16] = -8'd24;
        rom[62][17] = 8'd7;
        rom[62][18] = 8'd27;
        rom[62][19] = -8'd49;
        rom[62][20] = 8'd1;
        rom[62][21] = 8'd10;
        rom[62][22] = -8'd95;
        rom[62][23] = -8'd12;
        rom[62][24] = -8'd12;
        rom[62][25] = 8'd39;
        rom[62][26] = -8'd65;
        rom[62][27] = -8'd51;
        rom[62][28] = -8'd6;
        rom[62][29] = -8'd30;
        rom[62][30] = 8'd38;
        rom[62][31] = -8'd35;
        rom[62][32] = 8'd6;
        rom[62][33] = -8'd40;
        rom[62][34] = 8'd20;
        rom[62][35] = -8'd18;
        rom[62][36] = 8'd19;
        rom[62][37] = -8'd22;
        rom[62][38] = -8'd18;
        rom[62][39] = -8'd13;
        rom[62][40] = -8'd2;
        rom[62][41] = 8'd6;
        rom[62][42] = -8'd57;
        rom[62][43] = -8'd41;
        rom[62][44] = -8'd6;
        rom[62][45] = -8'd2;
        rom[62][46] = 8'd0;
        rom[62][47] = -8'd30;
        rom[62][48] = -8'd5;
        rom[62][49] = -8'd6;
        rom[62][50] = 8'd23;
        rom[62][51] = 8'd18;
        rom[62][52] = 8'd30;
        rom[62][53] = 8'd1;
        rom[62][54] = 8'd0;
        rom[62][55] = -8'd8;
        rom[62][56] = -8'd32;
        rom[62][57] = -8'd23;
        rom[62][58] = -8'd60;
        rom[62][59] = -8'd5;
        rom[62][60] = -8'd5;
        rom[62][61] = 8'd2;
        rom[62][62] = 8'd10;
        rom[62][63] = -8'd19;
        rom[63][0] = -8'd31;
        rom[63][1] = -8'd32;
        rom[63][2] = 8'd4;
        rom[63][3] = 8'd3;
        rom[63][4] = 8'd19;
        rom[63][5] = 8'd12;
        rom[63][6] = 8'd10;
        rom[63][7] = -8'd5;
        rom[63][8] = -8'd26;
        rom[63][9] = 8'd6;
        rom[63][10] = -8'd13;
        rom[63][11] = -8'd6;
        rom[63][12] = 8'd7;
        rom[63][13] = -8'd11;
        rom[63][14] = -8'd9;
        rom[63][15] = -8'd9;
        rom[63][16] = -8'd6;
        rom[63][17] = -8'd42;
        rom[63][18] = 8'd1;
        rom[63][19] = -8'd43;
        rom[63][20] = -8'd12;
        rom[63][21] = 8'd20;
        rom[63][22] = -8'd74;
        rom[63][23] = 8'd1;
        rom[63][24] = 8'd39;
        rom[63][25] = -8'd25;
        rom[63][26] = -8'd5;
        rom[63][27] = -8'd35;
        rom[63][28] = -8'd15;
        rom[63][29] = -8'd48;
        rom[63][30] = -8'd13;
        rom[63][31] = -8'd10;
        rom[63][32] = -8'd20;
        rom[63][33] = -8'd59;
        rom[63][34] = -8'd51;
        rom[63][35] = -8'd7;
        rom[63][36] = -8'd27;
        rom[63][37] = -8'd6;
        rom[63][38] = 8'd3;
        rom[63][39] = 8'd39;
        rom[63][40] = 8'd0;
        rom[63][41] = 8'd21;
        rom[63][42] = -8'd15;
        rom[63][43] = 8'd13;
        rom[63][44] = -8'd24;
        rom[63][45] = 8'd38;
        rom[63][46] = 8'd32;
        rom[63][47] = 8'd4;
        rom[63][48] = -8'd16;
        rom[63][49] = 8'd26;
        rom[63][50] = -8'd44;
        rom[63][51] = -8'd8;
        rom[63][52] = -8'd10;
        rom[63][53] = -8'd15;
        rom[63][54] = -8'd53;
        rom[63][55] = -8'd51;
        rom[63][56] = 8'd7;
        rom[63][57] = -8'd16;
        rom[63][58] = -8'd17;
        rom[63][59] = -8'd4;
        rom[63][60] = -8'd32;
        rom[63][61] = -8'd9;
        rom[63][62] = 8'd2;
        rom[63][63] = 8'd15;
        rom[64][0] = -8'd14;
        rom[64][1] = 8'd35;
        rom[64][2] = -8'd3;
        rom[64][3] = -8'd65;
        rom[64][4] = -8'd18;
        rom[64][5] = -8'd28;
        rom[64][6] = -8'd44;
        rom[64][7] = 8'd8;
        rom[64][8] = 8'd29;
        rom[64][9] = -8'd19;
        rom[64][10] = 8'd27;
        rom[64][11] = -8'd12;
        rom[64][12] = 8'd12;
        rom[64][13] = -8'd13;
        rom[64][14] = -8'd7;
        rom[64][15] = -8'd12;
        rom[64][16] = 8'd4;
        rom[64][17] = -8'd8;
        rom[64][18] = -8'd2;
        rom[64][19] = -8'd10;
        rom[64][20] = -8'd11;
        rom[64][21] = -8'd40;
        rom[64][22] = -8'd23;
        rom[64][23] = -8'd46;
        rom[64][24] = 8'd35;
        rom[64][25] = -8'd16;
        rom[64][26] = -8'd3;
        rom[64][27] = -8'd58;
        rom[64][28] = -8'd5;
        rom[64][29] = 8'd16;
        rom[64][30] = 8'd1;
        rom[64][31] = -8'd8;
        rom[64][32] = -8'd1;
        rom[64][33] = -8'd37;
        rom[64][34] = -8'd10;
        rom[64][35] = -8'd2;
        rom[64][36] = -8'd31;
        rom[64][37] = -8'd3;
        rom[64][38] = 8'd4;
        rom[64][39] = 8'd16;
        rom[64][40] = 8'd31;
        rom[64][41] = -8'd4;
        rom[64][42] = -8'd19;
        rom[64][43] = -8'd22;
        rom[64][44] = -8'd14;
        rom[64][45] = -8'd2;
        rom[64][46] = -8'd33;
        rom[64][47] = 8'd13;
        rom[64][48] = -8'd51;
        rom[64][49] = 8'd21;
        rom[64][50] = -8'd37;
        rom[64][51] = -8'd12;
        rom[64][52] = 8'd7;
        rom[64][53] = -8'd2;
        rom[64][54] = -8'd33;
        rom[64][55] = -8'd4;
        rom[64][56] = -8'd12;
        rom[64][57] = 8'd25;
        rom[64][58] = 8'd1;
        rom[64][59] = -8'd24;
        rom[64][60] = -8'd28;
        rom[64][61] = 8'd57;
        rom[64][62] = -8'd19;
        rom[64][63] = 8'd10;
        rom[65][0] = -8'd28;
        rom[65][1] = 8'd6;
        rom[65][2] = 8'd12;
        rom[65][3] = -8'd36;
        rom[65][4] = 8'd28;
        rom[65][5] = -8'd65;
        rom[65][6] = -8'd17;
        rom[65][7] = -8'd74;
        rom[65][8] = 8'd21;
        rom[65][9] = -8'd3;
        rom[65][10] = -8'd60;
        rom[65][11] = 8'd6;
        rom[65][12] = -8'd30;
        rom[65][13] = -8'd19;
        rom[65][14] = 8'd10;
        rom[65][15] = -8'd20;
        rom[65][16] = -8'd4;
        rom[65][17] = -8'd3;
        rom[65][18] = -8'd27;
        rom[65][19] = -8'd25;
        rom[65][20] = -8'd16;
        rom[65][21] = 8'd14;
        rom[65][22] = -8'd54;
        rom[65][23] = -8'd40;
        rom[65][24] = -8'd19;
        rom[65][25] = 8'd6;
        rom[65][26] = 8'd8;
        rom[65][27] = -8'd69;
        rom[65][28] = -8'd47;
        rom[65][29] = 8'd39;
        rom[65][30] = 8'd5;
        rom[65][31] = -8'd23;
        rom[65][32] = -8'd50;
        rom[65][33] = -8'd18;
        rom[65][34] = -8'd14;
        rom[65][35] = -8'd8;
        rom[65][36] = -8'd19;
        rom[65][37] = -8'd11;
        rom[65][38] = -8'd34;
        rom[65][39] = -8'd7;
        rom[65][40] = -8'd29;
        rom[65][41] = -8'd23;
        rom[65][42] = -8'd5;
        rom[65][43] = -8'd19;
        rom[65][44] = -8'd39;
        rom[65][45] = -8'd73;
        rom[65][46] = 8'd6;
        rom[65][47] = 8'd15;
        rom[65][48] = -8'd55;
        rom[65][49] = -8'd8;
        rom[65][50] = 8'd3;
        rom[65][51] = 8'd25;
        rom[65][52] = -8'd12;
        rom[65][53] = -8'd21;
        rom[65][54] = 8'd25;
        rom[65][55] = -8'd40;
        rom[65][56] = 8'd27;
        rom[65][57] = 8'd17;
        rom[65][58] = -8'd8;
        rom[65][59] = -8'd22;
        rom[65][60] = -8'd20;
        rom[65][61] = -8'd23;
        rom[65][62] = 8'd8;
        rom[65][63] = 8'd8;
        rom[66][0] = -8'd25;
        rom[66][1] = -8'd25;
        rom[66][2] = 8'd2;
        rom[66][3] = -8'd30;
        rom[66][4] = 8'd4;
        rom[66][5] = -8'd63;
        rom[66][6] = 8'd5;
        rom[66][7] = -8'd1;
        rom[66][8] = 8'd18;
        rom[66][9] = 8'd24;
        rom[66][10] = 8'd12;
        rom[66][11] = -8'd29;
        rom[66][12] = -8'd69;
        rom[66][13] = -8'd7;
        rom[66][14] = -8'd11;
        rom[66][15] = 8'd4;
        rom[66][16] = -8'd29;
        rom[66][17] = -8'd23;
        rom[66][18] = -8'd5;
        rom[66][19] = -8'd20;
        rom[66][20] = -8'd6;
        rom[66][21] = -8'd37;
        rom[66][22] = -8'd20;
        rom[66][23] = -8'd14;
        rom[66][24] = 8'd9;
        rom[66][25] = 8'd1;
        rom[66][26] = -8'd10;
        rom[66][27] = -8'd26;
        rom[66][28] = -8'd1;
        rom[66][29] = 8'd12;
        rom[66][30] = 8'd28;
        rom[66][31] = -8'd1;
        rom[66][32] = -8'd50;
        rom[66][33] = -8'd14;
        rom[66][34] = 8'd10;
        rom[66][35] = -8'd76;
        rom[66][36] = 8'd22;
        rom[66][37] = 8'd6;
        rom[66][38] = 8'd11;
        rom[66][39] = 8'd6;
        rom[66][40] = -8'd18;
        rom[66][41] = 8'd6;
        rom[66][42] = -8'd8;
        rom[66][43] = -8'd46;
        rom[66][44] = -8'd103;
        rom[66][45] = 8'd1;
        rom[66][46] = -8'd42;
        rom[66][47] = 8'd5;
        rom[66][48] = 8'd25;
        rom[66][49] = -8'd3;
        rom[66][50] = 8'd4;
        rom[66][51] = 8'd20;
        rom[66][52] = 8'd34;
        rom[66][53] = -8'd17;
        rom[66][54] = 8'd4;
        rom[66][55] = 8'd29;
        rom[66][56] = 8'd6;
        rom[66][57] = 8'd13;
        rom[66][58] = 8'd11;
        rom[66][59] = -8'd33;
        rom[66][60] = -8'd26;
        rom[66][61] = 8'd30;
        rom[66][62] = 8'd27;
        rom[66][63] = -8'd20;
        rom[67][0] = -8'd17;
        rom[67][1] = -8'd2;
        rom[67][2] = 8'd16;
        rom[67][3] = 8'd6;
        rom[67][4] = -8'd1;
        rom[67][5] = 8'd11;
        rom[67][6] = 8'd39;
        rom[67][7] = -8'd11;
        rom[67][8] = -8'd45;
        rom[67][9] = -8'd30;
        rom[67][10] = 8'd20;
        rom[67][11] = 8'd20;
        rom[67][12] = 8'd28;
        rom[67][13] = 8'd29;
        rom[67][14] = -8'd4;
        rom[67][15] = 8'd22;
        rom[67][16] = 8'd27;
        rom[67][17] = -8'd62;
        rom[67][18] = 8'd38;
        rom[67][19] = 8'd54;
        rom[67][20] = -8'd4;
        rom[67][21] = -8'd32;
        rom[67][22] = -8'd3;
        rom[67][23] = -8'd5;
        rom[67][24] = 8'd13;
        rom[67][25] = 8'd2;
        rom[67][26] = -8'd27;
        rom[67][27] = -8'd13;
        rom[67][28] = 8'd7;
        rom[67][29] = 8'd4;
        rom[67][30] = -8'd8;
        rom[67][31] = -8'd21;
        rom[67][32] = 8'd13;
        rom[67][33] = -8'd8;
        rom[67][34] = -8'd63;
        rom[67][35] = 8'd17;
        rom[67][36] = -8'd22;
        rom[67][37] = 8'd0;
        rom[67][38] = 8'd25;
        rom[67][39] = 8'd7;
        rom[67][40] = -8'd4;
        rom[67][41] = 8'd28;
        rom[67][42] = -8'd27;
        rom[67][43] = 8'd12;
        rom[67][44] = 8'd26;
        rom[67][45] = -8'd11;
        rom[67][46] = 8'd13;
        rom[67][47] = 8'd35;
        rom[67][48] = -8'd7;
        rom[67][49] = 8'd21;
        rom[67][50] = 8'd20;
        rom[67][51] = -8'd15;
        rom[67][52] = -8'd2;
        rom[67][53] = -8'd13;
        rom[67][54] = 8'd9;
        rom[67][55] = -8'd22;
        rom[67][56] = 8'd12;
        rom[67][57] = -8'd45;
        rom[67][58] = 8'd20;
        rom[67][59] = -8'd7;
        rom[67][60] = -8'd5;
        rom[67][61] = 8'd1;
        rom[67][62] = -8'd7;
        rom[67][63] = 8'd23;
        rom[68][0] = -8'd2;
        rom[68][1] = -8'd12;
        rom[68][2] = 8'd20;
        rom[68][3] = 8'd11;
        rom[68][4] = 8'd6;
        rom[68][5] = 8'd18;
        rom[68][6] = -8'd6;
        rom[68][7] = -8'd18;
        rom[68][8] = 8'd18;
        rom[68][9] = 8'd14;
        rom[68][10] = -8'd33;
        rom[68][11] = 8'd41;
        rom[68][12] = -8'd17;
        rom[68][13] = -8'd29;
        rom[68][14] = 8'd27;
        rom[68][15] = -8'd23;
        rom[68][16] = 8'd20;
        rom[68][17] = 8'd26;
        rom[68][18] = -8'd55;
        rom[68][19] = 8'd19;
        rom[68][20] = -8'd11;
        rom[68][21] = -8'd29;
        rom[68][22] = 8'd17;
        rom[68][23] = 8'd0;
        rom[68][24] = -8'd10;
        rom[68][25] = 8'd7;
        rom[68][26] = 8'd10;
        rom[68][27] = 8'd2;
        rom[68][28] = -8'd5;
        rom[68][29] = -8'd21;
        rom[68][30] = -8'd46;
        rom[68][31] = -8'd2;
        rom[68][32] = -8'd1;
        rom[68][33] = -8'd11;
        rom[68][34] = -8'd12;
        rom[68][35] = 8'd2;
        rom[68][36] = -8'd49;
        rom[68][37] = -8'd24;
        rom[68][38] = -8'd26;
        rom[68][39] = 8'd5;
        rom[68][40] = 8'd4;
        rom[68][41] = 8'd13;
        rom[68][42] = 8'd6;
        rom[68][43] = -8'd1;
        rom[68][44] = -8'd8;
        rom[68][45] = -8'd33;
        rom[68][46] = -8'd14;
        rom[68][47] = -8'd60;
        rom[68][48] = -8'd2;
        rom[68][49] = 8'd9;
        rom[68][50] = 8'd6;
        rom[68][51] = -8'd5;
        rom[68][52] = -8'd36;
        rom[68][53] = 8'd8;
        rom[68][54] = -8'd26;
        rom[68][55] = 8'd25;
        rom[68][56] = -8'd44;
        rom[68][57] = 8'd3;
        rom[68][58] = -8'd19;
        rom[68][59] = 8'd9;
        rom[68][60] = 8'd5;
        rom[68][61] = 8'd16;
        rom[68][62] = -8'd36;
        rom[68][63] = -8'd13;
        rom[69][0] = 8'd1;
        rom[69][1] = 8'd1;
        rom[69][2] = 8'd5;
        rom[69][3] = -8'd5;
        rom[69][4] = 8'd0;
        rom[69][5] = 8'd11;
        rom[69][6] = -8'd3;
        rom[69][7] = 8'd9;
        rom[69][8] = 8'd4;
        rom[69][9] = -8'd2;
        rom[69][10] = -8'd7;
        rom[69][11] = 8'd6;
        rom[69][12] = 8'd0;
        rom[69][13] = 8'd0;
        rom[69][14] = 8'd12;
        rom[69][15] = -8'd5;
        rom[69][16] = 8'd7;
        rom[69][17] = 8'd2;
        rom[69][18] = 8'd1;
        rom[69][19] = 8'd4;
        rom[69][20] = 8'd1;
        rom[69][21] = 8'd1;
        rom[69][22] = 8'd7;
        rom[69][23] = 8'd6;
        rom[69][24] = -8'd2;
        rom[69][25] = -8'd6;
        rom[69][26] = -8'd8;
        rom[69][27] = -8'd5;
        rom[69][28] = -8'd6;
        rom[69][29] = 8'd4;
        rom[69][30] = 8'd2;
        rom[69][31] = 8'd9;
        rom[69][32] = 8'd9;
        rom[69][33] = 8'd5;
        rom[69][34] = 8'd2;
        rom[69][35] = 8'd7;
        rom[69][36] = 8'd5;
        rom[69][37] = -8'd15;
        rom[69][38] = -8'd8;
        rom[69][39] = 8'd1;
        rom[69][40] = -8'd10;
        rom[69][41] = -8'd4;
        rom[69][42] = 8'd0;
        rom[69][43] = -8'd7;
        rom[69][44] = -8'd3;
        rom[69][45] = 8'd4;
        rom[69][46] = 8'd7;
        rom[69][47] = -8'd2;
        rom[69][48] = -8'd9;
        rom[69][49] = 8'd1;
        rom[69][50] = -8'd8;
        rom[69][51] = 8'd0;
        rom[69][52] = 8'd4;
        rom[69][53] = 8'd6;
        rom[69][54] = -8'd1;
        rom[69][55] = -8'd11;
        rom[69][56] = 8'd4;
        rom[69][57] = -8'd4;
        rom[69][58] = 8'd4;
        rom[69][59] = 8'd6;
        rom[69][60] = -8'd4;
        rom[69][61] = -8'd3;
        rom[69][62] = -8'd2;
        rom[69][63] = 8'd5;
        rom[70][0] = 8'd11;
        rom[70][1] = 8'd13;
        rom[70][2] = 8'd19;
        rom[70][3] = 8'd27;
        rom[70][4] = -8'd10;
        rom[70][5] = 8'd12;
        rom[70][6] = 8'd5;
        rom[70][7] = -8'd30;
        rom[70][8] = 8'd24;
        rom[70][9] = 8'd1;
        rom[70][10] = -8'd55;
        rom[70][11] = -8'd12;
        rom[70][12] = -8'd25;
        rom[70][13] = -8'd29;
        rom[70][14] = 8'd29;
        rom[70][15] = -8'd22;
        rom[70][16] = 8'd33;
        rom[70][17] = -8'd45;
        rom[70][18] = 8'd15;
        rom[70][19] = 8'd11;
        rom[70][20] = -8'd2;
        rom[70][21] = -8'd15;
        rom[70][22] = 8'd1;
        rom[70][23] = 8'd18;
        rom[70][24] = -8'd11;
        rom[70][25] = -8'd42;
        rom[70][26] = 8'd21;
        rom[70][27] = -8'd16;
        rom[70][28] = -8'd7;
        rom[70][29] = 8'd4;
        rom[70][30] = -8'd4;
        rom[70][31] = -8'd9;
        rom[70][32] = 8'd13;
        rom[70][33] = 8'd13;
        rom[70][34] = 8'd12;
        rom[70][35] = -8'd2;
        rom[70][36] = 8'd1;
        rom[70][37] = -8'd36;
        rom[70][38] = 8'd8;
        rom[70][39] = -8'd19;
        rom[70][40] = -8'd33;
        rom[70][41] = 8'd1;
        rom[70][42] = 8'd47;
        rom[70][43] = -8'd22;
        rom[70][44] = 8'd1;
        rom[70][45] = -8'd9;
        rom[70][46] = -8'd36;
        rom[70][47] = -8'd43;
        rom[70][48] = 8'd11;
        rom[70][49] = 8'd5;
        rom[70][50] = 8'd22;
        rom[70][51] = 8'd19;
        rom[70][52] = -8'd41;
        rom[70][53] = -8'd7;
        rom[70][54] = 8'd5;
        rom[70][55] = -8'd40;
        rom[70][56] = -8'd2;
        rom[70][57] = -8'd5;
        rom[70][58] = -8'd2;
        rom[70][59] = -8'd58;
        rom[70][60] = -8'd1;
        rom[70][61] = 8'd4;
        rom[70][62] = -8'd14;
        rom[70][63] = -8'd9;
        rom[71][0] = -8'd17;
        rom[71][1] = 8'd10;
        rom[71][2] = -8'd59;
        rom[71][3] = 8'd34;
        rom[71][4] = 8'd13;
        rom[71][5] = -8'd11;
        rom[71][6] = -8'd3;
        rom[71][7] = -8'd27;
        rom[71][8] = -8'd19;
        rom[71][9] = 8'd46;
        rom[71][10] = -8'd2;
        rom[71][11] = -8'd39;
        rom[71][12] = 8'd2;
        rom[71][13] = -8'd6;
        rom[71][14] = -8'd28;
        rom[71][15] = -8'd34;
        rom[71][16] = 8'd18;
        rom[71][17] = 8'd19;
        rom[71][18] = -8'd31;
        rom[71][19] = 8'd7;
        rom[71][20] = -8'd2;
        rom[71][21] = 8'd58;
        rom[71][22] = 8'd22;
        rom[71][23] = -8'd25;
        rom[71][24] = 8'd10;
        rom[71][25] = -8'd13;
        rom[71][26] = 8'd17;
        rom[71][27] = -8'd46;
        rom[71][28] = 8'd19;
        rom[71][29] = -8'd9;
        rom[71][30] = -8'd4;
        rom[71][31] = 8'd7;
        rom[71][32] = 8'd6;
        rom[71][33] = -8'd8;
        rom[71][34] = -8'd28;
        rom[71][35] = -8'd66;
        rom[71][36] = -8'd20;
        rom[71][37] = 8'd23;
        rom[71][38] = 8'd34;
        rom[71][39] = -8'd25;
        rom[71][40] = 8'd8;
        rom[71][41] = -8'd68;
        rom[71][42] = 8'd5;
        rom[71][43] = 8'd11;
        rom[71][44] = 8'd43;
        rom[71][45] = 8'd0;
        rom[71][46] = 8'd33;
        rom[71][47] = 8'd9;
        rom[71][48] = 8'd26;
        rom[71][49] = 8'd5;
        rom[71][50] = -8'd7;
        rom[71][51] = -8'd19;
        rom[71][52] = 8'd11;
        rom[71][53] = -8'd29;
        rom[71][54] = -8'd46;
        rom[71][55] = 8'd16;
        rom[71][56] = -8'd12;
        rom[71][57] = 8'd6;
        rom[71][58] = -8'd20;
        rom[71][59] = -8'd9;
        rom[71][60] = -8'd12;
        rom[71][61] = -8'd64;
        rom[71][62] = 8'd22;
        rom[71][63] = -8'd6;
        rom[72][0] = 8'd23;
        rom[72][1] = 8'd41;
        rom[72][2] = 8'd2;
        rom[72][3] = 8'd35;
        rom[72][4] = -8'd5;
        rom[72][5] = -8'd9;
        rom[72][6] = -8'd2;
        rom[72][7] = 8'd28;
        rom[72][8] = -8'd5;
        rom[72][9] = 8'd10;
        rom[72][10] = -8'd8;
        rom[72][11] = -8'd51;
        rom[72][12] = 8'd15;
        rom[72][13] = -8'd9;
        rom[72][14] = 8'd7;
        rom[72][15] = 8'd48;
        rom[72][16] = 8'd8;
        rom[72][17] = 8'd33;
        rom[72][18] = -8'd63;
        rom[72][19] = 8'd19;
        rom[72][20] = -8'd1;
        rom[72][21] = -8'd12;
        rom[72][22] = 8'd16;
        rom[72][23] = 8'd11;
        rom[72][24] = -8'd15;
        rom[72][25] = 8'd26;
        rom[72][26] = 8'd4;
        rom[72][27] = -8'd14;
        rom[72][28] = -8'd7;
        rom[72][29] = -8'd14;
        rom[72][30] = -8'd10;
        rom[72][31] = 8'd20;
        rom[72][32] = 8'd13;
        rom[72][33] = -8'd1;
        rom[72][34] = -8'd36;
        rom[72][35] = -8'd4;
        rom[72][36] = -8'd9;
        rom[72][37] = 8'd24;
        rom[72][38] = -8'd11;
        rom[72][39] = -8'd34;
        rom[72][40] = -8'd8;
        rom[72][41] = 8'd23;
        rom[72][42] = 8'd31;
        rom[72][43] = 8'd11;
        rom[72][44] = -8'd11;
        rom[72][45] = 8'd1;
        rom[72][46] = 8'd33;
        rom[72][47] = -8'd9;
        rom[72][48] = -8'd1;
        rom[72][49] = -8'd76;
        rom[72][50] = 8'd9;
        rom[72][51] = -8'd3;
        rom[72][52] = -8'd14;
        rom[72][53] = -8'd53;
        rom[72][54] = -8'd18;
        rom[72][55] = 8'd0;
        rom[72][56] = 8'd11;
        rom[72][57] = -8'd39;
        rom[72][58] = 8'd4;
        rom[72][59] = -8'd11;
        rom[72][60] = -8'd9;
        rom[72][61] = -8'd89;
        rom[72][62] = -8'd27;
        rom[72][63] = -8'd40;
        rom[73][0] = 8'd10;
        rom[73][1] = 8'd14;
        rom[73][2] = -8'd35;
        rom[73][3] = 8'd9;
        rom[73][4] = -8'd16;
        rom[73][5] = -8'd2;
        rom[73][6] = -8'd9;
        rom[73][7] = -8'd5;
        rom[73][8] = -8'd61;
        rom[73][9] = 8'd18;
        rom[73][10] = -8'd24;
        rom[73][11] = 8'd7;
        rom[73][12] = 8'd20;
        rom[73][13] = -8'd6;
        rom[73][14] = 8'd32;
        rom[73][15] = 8'd1;
        rom[73][16] = 8'd32;
        rom[73][17] = 8'd20;
        rom[73][18] = 8'd25;
        rom[73][19] = 8'd8;
        rom[73][20] = -8'd5;
        rom[73][21] = 8'd22;
        rom[73][22] = 8'd0;
        rom[73][23] = -8'd3;
        rom[73][24] = 8'd17;
        rom[73][25] = -8'd43;
        rom[73][26] = 8'd8;
        rom[73][27] = 8'd2;
        rom[73][28] = -8'd41;
        rom[73][29] = 8'd47;
        rom[73][30] = -8'd2;
        rom[73][31] = 8'd27;
        rom[73][32] = 8'd16;
        rom[73][33] = -8'd17;
        rom[73][34] = -8'd6;
        rom[73][35] = -8'd27;
        rom[73][36] = -8'd38;
        rom[73][37] = 8'd26;
        rom[73][38] = 8'd16;
        rom[73][39] = -8'd24;
        rom[73][40] = -8'd5;
        rom[73][41] = -8'd12;
        rom[73][42] = 8'd36;
        rom[73][43] = 8'd4;
        rom[73][44] = -8'd23;
        rom[73][45] = 8'd26;
        rom[73][46] = -8'd26;
        rom[73][47] = -8'd23;
        rom[73][48] = -8'd5;
        rom[73][49] = -8'd4;
        rom[73][50] = -8'd84;
        rom[73][51] = -8'd43;
        rom[73][52] = 8'd2;
        rom[73][53] = 8'd19;
        rom[73][54] = -8'd50;
        rom[73][55] = 8'd25;
        rom[73][56] = -8'd14;
        rom[73][57] = -8'd33;
        rom[73][58] = -8'd35;
        rom[73][59] = 8'd5;
        rom[73][60] = 8'd17;
        rom[73][61] = -8'd2;
        rom[73][62] = 8'd4;
        rom[73][63] = -8'd39;
        rom[74][0] = -8'd19;
        rom[74][1] = 8'd19;
        rom[74][2] = 8'd13;
        rom[74][3] = 8'd10;
        rom[74][4] = -8'd16;
        rom[74][5] = -8'd10;
        rom[74][6] = 8'd44;
        rom[74][7] = -8'd32;
        rom[74][8] = 8'd13;
        rom[74][9] = -8'd22;
        rom[74][10] = 8'd33;
        rom[74][11] = -8'd1;
        rom[74][12] = 8'd14;
        rom[74][13] = -8'd55;
        rom[74][14] = 8'd5;
        rom[74][15] = -8'd5;
        rom[74][16] = -8'd25;
        rom[74][17] = -8'd30;
        rom[74][18] = 8'd4;
        rom[74][19] = -8'd14;
        rom[74][20] = -8'd7;
        rom[74][21] = 8'd13;
        rom[74][22] = -8'd30;
        rom[74][23] = -8'd49;
        rom[74][24] = 8'd16;
        rom[74][25] = 8'd12;
        rom[74][26] = -8'd8;
        rom[74][27] = -8'd34;
        rom[74][28] = -8'd20;
        rom[74][29] = -8'd17;
        rom[74][30] = 8'd11;
        rom[74][31] = -8'd16;
        rom[74][32] = -8'd15;
        rom[74][33] = 8'd5;
        rom[74][34] = -8'd32;
        rom[74][35] = -8'd21;
        rom[74][36] = 8'd33;
        rom[74][37] = -8'd59;
        rom[74][38] = 8'd16;
        rom[74][39] = 8'd36;
        rom[74][40] = -8'd6;
        rom[74][41] = -8'd22;
        rom[74][42] = -8'd21;
        rom[74][43] = -8'd37;
        rom[74][44] = 8'd0;
        rom[74][45] = -8'd24;
        rom[74][46] = 8'd11;
        rom[74][47] = 8'd7;
        rom[74][48] = 8'd23;
        rom[74][49] = 8'd20;
        rom[74][50] = -8'd9;
        rom[74][51] = -8'd5;
        rom[74][52] = -8'd5;
        rom[74][53] = -8'd44;
        rom[74][54] = -8'd17;
        rom[74][55] = -8'd34;
        rom[74][56] = -8'd33;
        rom[74][57] = 8'd20;
        rom[74][58] = 8'd9;
        rom[74][59] = -8'd36;
        rom[74][60] = 8'd17;
        rom[74][61] = 8'd2;
        rom[74][62] = 8'd3;
        rom[74][63] = 8'd8;
        rom[75][0] = 8'd26;
        rom[75][1] = 8'd11;
        rom[75][2] = 8'd13;
        rom[75][3] = -8'd34;
        rom[75][4] = 8'd8;
        rom[75][5] = 8'd18;
        rom[75][6] = -8'd13;
        rom[75][7] = 8'd6;
        rom[75][8] = -8'd23;
        rom[75][9] = -8'd27;
        rom[75][10] = -8'd4;
        rom[75][11] = -8'd32;
        rom[75][12] = 8'd31;
        rom[75][13] = 8'd16;
        rom[75][14] = 8'd24;
        rom[75][15] = -8'd2;
        rom[75][16] = -8'd43;
        rom[75][17] = -8'd71;
        rom[75][18] = 8'd10;
        rom[75][19] = 8'd32;
        rom[75][20] = -8'd4;
        rom[75][21] = 8'd6;
        rom[75][22] = 8'd41;
        rom[75][23] = -8'd1;
        rom[75][24] = 8'd14;
        rom[75][25] = -8'd65;
        rom[75][26] = 8'd37;
        rom[75][27] = 8'd37;
        rom[75][28] = 8'd13;
        rom[75][29] = 8'd43;
        rom[75][30] = -8'd43;
        rom[75][31] = 8'd38;
        rom[75][32] = -8'd53;
        rom[75][33] = -8'd10;
        rom[75][34] = 8'd29;
        rom[75][35] = 8'd27;
        rom[75][36] = 8'd35;
        rom[75][37] = -8'd1;
        rom[75][38] = -8'd18;
        rom[75][39] = 8'd8;
        rom[75][40] = 8'd3;
        rom[75][41] = -8'd12;
        rom[75][42] = 8'd45;
        rom[75][43] = 8'd24;
        rom[75][44] = 8'd27;
        rom[75][45] = 8'd14;
        rom[75][46] = 8'd36;
        rom[75][47] = 8'd31;
        rom[75][48] = 8'd22;
        rom[75][49] = -8'd16;
        rom[75][50] = -8'd21;
        rom[75][51] = 8'd11;
        rom[75][52] = -8'd14;
        rom[75][53] = -8'd19;
        rom[75][54] = 8'd19;
        rom[75][55] = -8'd7;
        rom[75][56] = 8'd25;
        rom[75][57] = 8'd20;
        rom[75][58] = 8'd23;
        rom[75][59] = 8'd4;
        rom[75][60] = -8'd35;
        rom[75][61] = 8'd4;
        rom[75][62] = 8'd43;
        rom[75][63] = 8'd21;
        rom[76][0] = 8'd19;
        rom[76][1] = -8'd40;
        rom[76][2] = 8'd39;
        rom[76][3] = -8'd38;
        rom[76][4] = -8'd15;
        rom[76][5] = 8'd7;
        rom[76][6] = 8'd5;
        rom[76][7] = -8'd26;
        rom[76][8] = -8'd16;
        rom[76][9] = 8'd22;
        rom[76][10] = 8'd24;
        rom[76][11] = -8'd14;
        rom[76][12] = -8'd53;
        rom[76][13] = 8'd44;
        rom[76][14] = -8'd4;
        rom[76][15] = -8'd44;
        rom[76][16] = -8'd27;
        rom[76][17] = -8'd20;
        rom[76][18] = 8'd2;
        rom[76][19] = -8'd90;
        rom[76][20] = -8'd7;
        rom[76][21] = -8'd20;
        rom[76][22] = -8'd27;
        rom[76][23] = -8'd5;
        rom[76][24] = -8'd23;
        rom[76][25] = 8'd16;
        rom[76][26] = -8'd9;
        rom[76][27] = -8'd2;
        rom[76][28] = 8'd21;
        rom[76][29] = -8'd3;
        rom[76][30] = 8'd8;
        rom[76][31] = 8'd22;
        rom[76][32] = -8'd23;
        rom[76][33] = -8'd80;
        rom[76][34] = -8'd2;
        rom[76][35] = -8'd55;
        rom[76][36] = 8'd19;
        rom[76][37] = -8'd1;
        rom[76][38] = 8'd9;
        rom[76][39] = 8'd5;
        rom[76][40] = 8'd25;
        rom[76][41] = 8'd0;
        rom[76][42] = -8'd10;
        rom[76][43] = -8'd6;
        rom[76][44] = 8'd6;
        rom[76][45] = -8'd72;
        rom[76][46] = -8'd41;
        rom[76][47] = -8'd1;
        rom[76][48] = 8'd28;
        rom[76][49] = 8'd27;
        rom[76][50] = 8'd34;
        rom[76][51] = 8'd13;
        rom[76][52] = -8'd24;
        rom[76][53] = -8'd45;
        rom[76][54] = -8'd32;
        rom[76][55] = 8'd9;
        rom[76][56] = 8'd1;
        rom[76][57] = 8'd34;
        rom[76][58] = 8'd4;
        rom[76][59] = -8'd37;
        rom[76][60] = -8'd20;
        rom[76][61] = 8'd3;
        rom[76][62] = 8'd12;
        rom[76][63] = 8'd21;
        rom[77][0] = 8'd19;
        rom[77][1] = -8'd25;
        rom[77][2] = 8'd14;
        rom[77][3] = -8'd51;
        rom[77][4] = 8'd20;
        rom[77][5] = -8'd12;
        rom[77][6] = -8'd34;
        rom[77][7] = 8'd1;
        rom[77][8] = 8'd8;
        rom[77][9] = -8'd36;
        rom[77][10] = 8'd9;
        rom[77][11] = -8'd7;
        rom[77][12] = -8'd2;
        rom[77][13] = 8'd20;
        rom[77][14] = 8'd24;
        rom[77][15] = 8'd0;
        rom[77][16] = -8'd20;
        rom[77][17] = -8'd44;
        rom[77][18] = 8'd13;
        rom[77][19] = -8'd6;
        rom[77][20] = 8'd2;
        rom[77][21] = 8'd9;
        rom[77][22] = -8'd30;
        rom[77][23] = 8'd23;
        rom[77][24] = -8'd9;
        rom[77][25] = -8'd42;
        rom[77][26] = -8'd13;
        rom[77][27] = 8'd13;
        rom[77][28] = -8'd2;
        rom[77][29] = 8'd9;
        rom[77][30] = -8'd12;
        rom[77][31] = -8'd2;
        rom[77][32] = 8'd1;
        rom[77][33] = -8'd25;
        rom[77][34] = -8'd58;
        rom[77][35] = -8'd8;
        rom[77][36] = -8'd43;
        rom[77][37] = -8'd26;
        rom[77][38] = -8'd21;
        rom[77][39] = 8'd41;
        rom[77][40] = -8'd15;
        rom[77][41] = 8'd2;
        rom[77][42] = -8'd13;
        rom[77][43] = 8'd16;
        rom[77][44] = 8'd0;
        rom[77][45] = 8'd15;
        rom[77][46] = 8'd13;
        rom[77][47] = -8'd25;
        rom[77][48] = 8'd0;
        rom[77][49] = -8'd40;
        rom[77][50] = -8'd45;
        rom[77][51] = 8'd13;
        rom[77][52] = 8'd19;
        rom[77][53] = -8'd25;
        rom[77][54] = 8'd5;
        rom[77][55] = 8'd1;
        rom[77][56] = -8'd8;
        rom[77][57] = 8'd12;
        rom[77][58] = -8'd8;
        rom[77][59] = -8'd20;
        rom[77][60] = -8'd36;
        rom[77][61] = 8'd26;
        rom[77][62] = -8'd35;
        rom[77][63] = 8'd25;
        rom[78][0] = 8'd32;
        rom[78][1] = 8'd22;
        rom[78][2] = 8'd0;
        rom[78][3] = 8'd31;
        rom[78][4] = -8'd18;
        rom[78][5] = -8'd28;
        rom[78][6] = -8'd13;
        rom[78][7] = -8'd27;
        rom[78][8] = -8'd8;
        rom[78][9] = -8'd37;
        rom[78][10] = 8'd17;
        rom[78][11] = -8'd19;
        rom[78][12] = 8'd21;
        rom[78][13] = -8'd7;
        rom[78][14] = 8'd6;
        rom[78][15] = 8'd16;
        rom[78][16] = 8'd9;
        rom[78][17] = -8'd43;
        rom[78][18] = -8'd56;
        rom[78][19] = 8'd10;
        rom[78][20] = -8'd4;
        rom[78][21] = -8'd22;
        rom[78][22] = -8'd15;
        rom[78][23] = -8'd3;
        rom[78][24] = -8'd40;
        rom[78][25] = 8'd9;
        rom[78][26] = 8'd2;
        rom[78][27] = -8'd6;
        rom[78][28] = -8'd48;
        rom[78][29] = -8'd65;
        rom[78][30] = -8'd28;
        rom[78][31] = 8'd6;
        rom[78][32] = 8'd14;
        rom[78][33] = 8'd30;
        rom[78][34] = -8'd14;
        rom[78][35] = 8'd21;
        rom[78][36] = -8'd33;
        rom[78][37] = 8'd8;
        rom[78][38] = -8'd50;
        rom[78][39] = 8'd26;
        rom[78][40] = 8'd48;
        rom[78][41] = 8'd0;
        rom[78][42] = 8'd3;
        rom[78][43] = -8'd9;
        rom[78][44] = -8'd18;
        rom[78][45] = 8'd35;
        rom[78][46] = 8'd22;
        rom[78][47] = -8'd30;
        rom[78][48] = -8'd4;
        rom[78][49] = -8'd12;
        rom[78][50] = 8'd15;
        rom[78][51] = -8'd18;
        rom[78][52] = -8'd6;
        rom[78][53] = 8'd3;
        rom[78][54] = 8'd9;
        rom[78][55] = -8'd77;
        rom[78][56] = 8'd24;
        rom[78][57] = 8'd1;
        rom[78][58] = -8'd22;
        rom[78][59] = 8'd7;
        rom[78][60] = -8'd33;
        rom[78][61] = 8'd2;
        rom[78][62] = 8'd13;
        rom[78][63] = -8'd12;
        rom[79][0] = -8'd3;
        rom[79][1] = -8'd46;
        rom[79][2] = -8'd34;
        rom[79][3] = -8'd24;
        rom[79][4] = -8'd31;
        rom[79][5] = 8'd1;
        rom[79][6] = 8'd4;
        rom[79][7] = -8'd10;
        rom[79][8] = -8'd67;
        rom[79][9] = -8'd19;
        rom[79][10] = -8'd74;
        rom[79][11] = -8'd13;
        rom[79][12] = 8'd54;
        rom[79][13] = 8'd24;
        rom[79][14] = -8'd4;
        rom[79][15] = -8'd13;
        rom[79][16] = -8'd12;
        rom[79][17] = 8'd30;
        rom[79][18] = 8'd14;
        rom[79][19] = 8'd4;
        rom[79][20] = 8'd6;
        rom[79][21] = -8'd11;
        rom[79][22] = -8'd32;
        rom[79][23] = 8'd10;
        rom[79][24] = 8'd9;
        rom[79][25] = 8'd6;
        rom[79][26] = -8'd5;
        rom[79][27] = -8'd27;
        rom[79][28] = -8'd12;
        rom[79][29] = 8'd3;
        rom[79][30] = -8'd16;
        rom[79][31] = -8'd22;
        rom[79][32] = 8'd28;
        rom[79][33] = 8'd31;
        rom[79][34] = -8'd10;
        rom[79][35] = 8'd11;
        rom[79][36] = 8'd19;
        rom[79][37] = -8'd1;
        rom[79][38] = 8'd1;
        rom[79][39] = 8'd0;
        rom[79][40] = -8'd16;
        rom[79][41] = 8'd12;
        rom[79][42] = 8'd3;
        rom[79][43] = -8'd42;
        rom[79][44] = -8'd23;
        rom[79][45] = -8'd45;
        rom[79][46] = 8'd34;
        rom[79][47] = -8'd3;
        rom[79][48] = -8'd16;
        rom[79][49] = -8'd14;
        rom[79][50] = -8'd22;
        rom[79][51] = -8'd35;
        rom[79][52] = 8'd9;
        rom[79][53] = -8'd4;
        rom[79][54] = 8'd29;
        rom[79][55] = 8'd15;
        rom[79][56] = 8'd11;
        rom[79][57] = 8'd6;
        rom[79][58] = -8'd18;
        rom[79][59] = -8'd26;
        rom[79][60] = -8'd35;
        rom[79][61] = -8'd21;
        rom[79][62] = -8'd7;
        rom[79][63] = -8'd10;
        rom[80][0] = 8'd4;
        rom[80][1] = -8'd1;
        rom[80][2] = -8'd2;
        rom[80][3] = -8'd4;
        rom[80][4] = -8'd1;
        rom[80][5] = 8'd8;
        rom[80][6] = 8'd6;
        rom[80][7] = 8'd8;
        rom[80][8] = -8'd9;
        rom[80][9] = 8'd0;
        rom[80][10] = -8'd6;
        rom[80][11] = 8'd6;
        rom[80][12] = 8'd3;
        rom[80][13] = 8'd4;
        rom[80][14] = 8'd1;
        rom[80][15] = 8'd7;
        rom[80][16] = 8'd3;
        rom[80][17] = -8'd4;
        rom[80][18] = -8'd3;
        rom[80][19] = -8'd7;
        rom[80][20] = 8'd0;
        rom[80][21] = -8'd5;
        rom[80][22] = -8'd4;
        rom[80][23] = 8'd7;
        rom[80][24] = -8'd6;
        rom[80][25] = 8'd1;
        rom[80][26] = -8'd3;
        rom[80][27] = -8'd5;
        rom[80][28] = -8'd5;
        rom[80][29] = 8'd9;
        rom[80][30] = 8'd2;
        rom[80][31] = 8'd4;
        rom[80][32] = 8'd4;
        rom[80][33] = 8'd3;
        rom[80][34] = 8'd9;
        rom[80][35] = 8'd6;
        rom[80][36] = -8'd1;
        rom[80][37] = -8'd6;
        rom[80][38] = 8'd4;
        rom[80][39] = 8'd0;
        rom[80][40] = -8'd2;
        rom[80][41] = 8'd7;
        rom[80][42] = -8'd2;
        rom[80][43] = 8'd9;
        rom[80][44] = 8'd6;
        rom[80][45] = 8'd7;
        rom[80][46] = -8'd2;
        rom[80][47] = -8'd4;
        rom[80][48] = -8'd3;
        rom[80][49] = -8'd5;
        rom[80][50] = -8'd6;
        rom[80][51] = -8'd5;
        rom[80][52] = -8'd9;
        rom[80][53] = -8'd6;
        rom[80][54] = 8'd7;
        rom[80][55] = -8'd9;
        rom[80][56] = 8'd3;
        rom[80][57] = -8'd1;
        rom[80][58] = -8'd1;
        rom[80][59] = -8'd2;
        rom[80][60] = 8'd4;
        rom[80][61] = 8'd5;
        rom[80][62] = 8'd5;
        rom[80][63] = -8'd5;
        rom[81][0] = 8'd46;
        rom[81][1] = 8'd18;
        rom[81][2] = 8'd38;
        rom[81][3] = 8'd48;
        rom[81][4] = 8'd26;
        rom[81][5] = 8'd38;
        rom[81][6] = 8'd49;
        rom[81][7] = 8'd49;
        rom[81][8] = 8'd18;
        rom[81][9] = -8'd28;
        rom[81][10] = -8'd81;
        rom[81][11] = -8'd3;
        rom[81][12] = 8'd14;
        rom[81][13] = -8'd21;
        rom[81][14] = 8'd24;
        rom[81][15] = 8'd45;
        rom[81][16] = 8'd43;
        rom[81][17] = 8'd14;
        rom[81][18] = 8'd15;
        rom[81][19] = 8'd10;
        rom[81][20] = -8'd2;
        rom[81][21] = -8'd37;
        rom[81][22] = 8'd41;
        rom[81][23] = 8'd30;
        rom[81][24] = 8'd20;
        rom[81][25] = 8'd9;
        rom[81][26] = -8'd36;
        rom[81][27] = 8'd5;
        rom[81][28] = -8'd23;
        rom[81][29] = -8'd15;
        rom[81][30] = 8'd8;
        rom[81][31] = 8'd23;
        rom[81][32] = 8'd25;
        rom[81][33] = -8'd15;
        rom[81][34] = 8'd10;
        rom[81][35] = 8'd2;
        rom[81][36] = 8'd30;
        rom[81][37] = 8'd21;
        rom[81][38] = 8'd1;
        rom[81][39] = 8'd11;
        rom[81][40] = 8'd38;
        rom[81][41] = 8'd23;
        rom[81][42] = 8'd1;
        rom[81][43] = 8'd7;
        rom[81][44] = -8'd9;
        rom[81][45] = -8'd4;
        rom[81][46] = -8'd25;
        rom[81][47] = -8'd42;
        rom[81][48] = 8'd15;
        rom[81][49] = 8'd4;
        rom[81][50] = -8'd2;
        rom[81][51] = -8'd44;
        rom[81][52] = -8'd1;
        rom[81][53] = 8'd38;
        rom[81][54] = -8'd5;
        rom[81][55] = 8'd0;
        rom[81][56] = -8'd30;
        rom[81][57] = -8'd24;
        rom[81][58] = -8'd60;
        rom[81][59] = 8'd2;
        rom[81][60] = -8'd28;
        rom[81][61] = 8'd64;
        rom[81][62] = -8'd84;
        rom[81][63] = -8'd25;
        rom[82][0] = 8'd10;
        rom[82][1] = -8'd4;
        rom[82][2] = 8'd2;
        rom[82][3] = 8'd39;
        rom[82][4] = -8'd34;
        rom[82][5] = 8'd12;
        rom[82][6] = -8'd21;
        rom[82][7] = 8'd32;
        rom[82][8] = -8'd29;
        rom[82][9] = 8'd13;
        rom[82][10] = -8'd1;
        rom[82][11] = 8'd9;
        rom[82][12] = 8'd5;
        rom[82][13] = 8'd10;
        rom[82][14] = -8'd5;
        rom[82][15] = -8'd14;
        rom[82][16] = 8'd9;
        rom[82][17] = 8'd5;
        rom[82][18] = 8'd19;
        rom[82][19] = -8'd20;
        rom[82][20] = -8'd13;
        rom[82][21] = -8'd9;
        rom[82][22] = 8'd19;
        rom[82][23] = -8'd1;
        rom[82][24] = 8'd23;
        rom[82][25] = 8'd5;
        rom[82][26] = -8'd30;
        rom[82][27] = 8'd24;
        rom[82][28] = -8'd5;
        rom[82][29] = -8'd14;
        rom[82][30] = 8'd1;
        rom[82][31] = 8'd16;
        rom[82][32] = -8'd48;
        rom[82][33] = 8'd8;
        rom[82][34] = -8'd5;
        rom[82][35] = 8'd11;
        rom[82][36] = -8'd20;
        rom[82][37] = 8'd14;
        rom[82][38] = -8'd1;
        rom[82][39] = 8'd31;
        rom[82][40] = 8'd1;
        rom[82][41] = 8'd25;
        rom[82][42] = -8'd8;
        rom[82][43] = -8'd21;
        rom[82][44] = -8'd20;
        rom[82][45] = 8'd19;
        rom[82][46] = -8'd34;
        rom[82][47] = 8'd3;
        rom[82][48] = -8'd20;
        rom[82][49] = -8'd6;
        rom[82][50] = 8'd11;
        rom[82][51] = -8'd6;
        rom[82][52] = -8'd4;
        rom[82][53] = -8'd29;
        rom[82][54] = -8'd12;
        rom[82][55] = -8'd53;
        rom[82][56] = 8'd12;
        rom[82][57] = -8'd46;
        rom[82][58] = -8'd33;
        rom[82][59] = 8'd18;
        rom[82][60] = -8'd6;
        rom[82][61] = -8'd23;
        rom[82][62] = -8'd17;
        rom[82][63] = -8'd11;
        rom[83][0] = -8'd43;
        rom[83][1] = -8'd6;
        rom[83][2] = -8'd69;
        rom[83][3] = -8'd59;
        rom[83][4] = -8'd22;
        rom[83][5] = 8'd23;
        rom[83][6] = 8'd19;
        rom[83][7] = 8'd10;
        rom[83][8] = -8'd24;
        rom[83][9] = 8'd8;
        rom[83][10] = -8'd17;
        rom[83][11] = -8'd19;
        rom[83][12] = -8'd11;
        rom[83][13] = -8'd69;
        rom[83][14] = 8'd2;
        rom[83][15] = 8'd3;
        rom[83][16] = 8'd10;
        rom[83][17] = 8'd9;
        rom[83][18] = 8'd13;
        rom[83][19] = -8'd9;
        rom[83][20] = 8'd3;
        rom[83][21] = 8'd25;
        rom[83][22] = -8'd46;
        rom[83][23] = -8'd29;
        rom[83][24] = -8'd6;
        rom[83][25] = 8'd10;
        rom[83][26] = -8'd6;
        rom[83][27] = -8'd62;
        rom[83][28] = 8'd64;
        rom[83][29] = -8'd7;
        rom[83][30] = 8'd19;
        rom[83][31] = -8'd3;
        rom[83][32] = -8'd9;
        rom[83][33] = -8'd33;
        rom[83][34] = -8'd4;
        rom[83][35] = 8'd10;
        rom[83][36] = -8'd28;
        rom[83][37] = -8'd13;
        rom[83][38] = -8'd20;
        rom[83][39] = -8'd27;
        rom[83][40] = -8'd9;
        rom[83][41] = -8'd18;
        rom[83][42] = -8'd63;
        rom[83][43] = -8'd4;
        rom[83][44] = 8'd14;
        rom[83][45] = -8'd48;
        rom[83][46] = -8'd7;
        rom[83][47] = 8'd18;
        rom[83][48] = -8'd4;
        rom[83][49] = -8'd37;
        rom[83][50] = -8'd70;
        rom[83][51] = -8'd17;
        rom[83][52] = 8'd10;
        rom[83][53] = 8'd3;
        rom[83][54] = 8'd20;
        rom[83][55] = 8'd14;
        rom[83][56] = 8'd27;
        rom[83][57] = 8'd16;
        rom[83][58] = 8'd32;
        rom[83][59] = 8'd4;
        rom[83][60] = 8'd7;
        rom[83][61] = 8'd11;
        rom[83][62] = -8'd5;
        rom[83][63] = 8'd1;
        rom[84][0] = -8'd7;
        rom[84][1] = -8'd6;
        rom[84][2] = 8'd10;
        rom[84][3] = 8'd26;
        rom[84][4] = 8'd34;
        rom[84][5] = -8'd5;
        rom[84][6] = -8'd13;
        rom[84][7] = -8'd60;
        rom[84][8] = 8'd11;
        rom[84][9] = 8'd15;
        rom[84][10] = -8'd26;
        rom[84][11] = -8'd17;
        rom[84][12] = -8'd76;
        rom[84][13] = -8'd17;
        rom[84][14] = 8'd1;
        rom[84][15] = -8'd28;
        rom[84][16] = -8'd22;
        rom[84][17] = -8'd24;
        rom[84][18] = -8'd58;
        rom[84][19] = -8'd3;
        rom[84][20] = 8'd3;
        rom[84][21] = 8'd2;
        rom[84][22] = 8'd7;
        rom[84][23] = 8'd16;
        rom[84][24] = -8'd5;
        rom[84][25] = -8'd37;
        rom[84][26] = 8'd20;
        rom[84][27] = 8'd2;
        rom[84][28] = -8'd4;
        rom[84][29] = 8'd16;
        rom[84][30] = -8'd6;
        rom[84][31] = -8'd3;
        rom[84][32] = -8'd27;
        rom[84][33] = -8'd36;
        rom[84][34] = -8'd12;
        rom[84][35] = 8'd5;
        rom[84][36] = -8'd28;
        rom[84][37] = 8'd2;
        rom[84][38] = -8'd9;
        rom[84][39] = -8'd30;
        rom[84][40] = 8'd1;
        rom[84][41] = -8'd47;
        rom[84][42] = 8'd8;
        rom[84][43] = 8'd1;
        rom[84][44] = -8'd20;
        rom[84][45] = -8'd4;
        rom[84][46] = -8'd34;
        rom[84][47] = 8'd40;
        rom[84][48] = -8'd10;
        rom[84][49] = -8'd10;
        rom[84][50] = 8'd21;
        rom[84][51] = -8'd12;
        rom[84][52] = -8'd5;
        rom[84][53] = 8'd6;
        rom[84][54] = -8'd13;
        rom[84][55] = -8'd5;
        rom[84][56] = 8'd2;
        rom[84][57] = -8'd24;
        rom[84][58] = 8'd30;
        rom[84][59] = -8'd26;
        rom[84][60] = 8'd11;
        rom[84][61] = -8'd14;
        rom[84][62] = 8'd34;
        rom[84][63] = -8'd11;
        rom[85][0] = 8'd8;
        rom[85][1] = -8'd8;
        rom[85][2] = 8'd5;
        rom[85][3] = 8'd3;
        rom[85][4] = 8'd7;
        rom[85][5] = 8'd9;
        rom[85][6] = 8'd6;
        rom[85][7] = -8'd5;
        rom[85][8] = -8'd4;
        rom[85][9] = -8'd6;
        rom[85][10] = 8'd8;
        rom[85][11] = -8'd5;
        rom[85][12] = 8'd2;
        rom[85][13] = 8'd8;
        rom[85][14] = 8'd0;
        rom[85][15] = -8'd8;
        rom[85][16] = -8'd1;
        rom[85][17] = -8'd4;
        rom[85][18] = -8'd2;
        rom[85][19] = 8'd5;
        rom[85][20] = -8'd3;
        rom[85][21] = -8'd8;
        rom[85][22] = -8'd6;
        rom[85][23] = 8'd1;
        rom[85][24] = 8'd1;
        rom[85][25] = 8'd3;
        rom[85][26] = -8'd7;
        rom[85][27] = 8'd8;
        rom[85][28] = -8'd11;
        rom[85][29] = -8'd1;
        rom[85][30] = 8'd5;
        rom[85][31] = -8'd1;
        rom[85][32] = -8'd9;
        rom[85][33] = 8'd1;
        rom[85][34] = -8'd1;
        rom[85][35] = 8'd9;
        rom[85][36] = -8'd1;
        rom[85][37] = 8'd9;
        rom[85][38] = 8'd3;
        rom[85][39] = -8'd8;
        rom[85][40] = -8'd7;
        rom[85][41] = -8'd3;
        rom[85][42] = -8'd8;
        rom[85][43] = -8'd3;
        rom[85][44] = -8'd4;
        rom[85][45] = 8'd8;
        rom[85][46] = 8'd2;
        rom[85][47] = 8'd8;
        rom[85][48] = 8'd1;
        rom[85][49] = -8'd6;
        rom[85][50] = -8'd2;
        rom[85][51] = -8'd1;
        rom[85][52] = -8'd4;
        rom[85][53] = -8'd1;
        rom[85][54] = -8'd5;
        rom[85][55] = 8'd7;
        rom[85][56] = -8'd8;
        rom[85][57] = 8'd7;
        rom[85][58] = 8'd0;
        rom[85][59] = -8'd3;
        rom[85][60] = 8'd9;
        rom[85][61] = 8'd5;
        rom[85][62] = 8'd5;
        rom[85][63] = 8'd2;
        rom[86][0] = -8'd14;
        rom[86][1] = 8'd11;
        rom[86][2] = -8'd25;
        rom[86][3] = -8'd7;
        rom[86][4] = 8'd0;
        rom[86][5] = -8'd35;
        rom[86][6] = -8'd35;
        rom[86][7] = 8'd13;
        rom[86][8] = 8'd6;
        rom[86][9] = -8'd15;
        rom[86][10] = 8'd36;
        rom[86][11] = -8'd32;
        rom[86][12] = -8'd7;
        rom[86][13] = -8'd6;
        rom[86][14] = 8'd5;
        rom[86][15] = -8'd22;
        rom[86][16] = -8'd55;
        rom[86][17] = -8'd28;
        rom[86][18] = -8'd66;
        rom[86][19] = 8'd30;
        rom[86][20] = -8'd2;
        rom[86][21] = -8'd11;
        rom[86][22] = -8'd8;
        rom[86][23] = -8'd26;
        rom[86][24] = -8'd1;
        rom[86][25] = -8'd1;
        rom[86][26] = 8'd7;
        rom[86][27] = -8'd8;
        rom[86][28] = 8'd11;
        rom[86][29] = 8'd0;
        rom[86][30] = -8'd19;
        rom[86][31] = -8'd10;
        rom[86][32] = -8'd5;
        rom[86][33] = -8'd11;
        rom[86][34] = 8'd14;
        rom[86][35] = -8'd13;
        rom[86][36] = 8'd7;
        rom[86][37] = -8'd13;
        rom[86][38] = -8'd40;
        rom[86][39] = -8'd16;
        rom[86][40] = -8'd21;
        rom[86][41] = 8'd21;
        rom[86][42] = -8'd7;
        rom[86][43] = 8'd32;
        rom[86][44] = -8'd7;
        rom[86][45] = -8'd21;
        rom[86][46] = 8'd29;
        rom[86][47] = -8'd20;
        rom[86][48] = -8'd52;
        rom[86][49] = -8'd25;
        rom[86][50] = 8'd28;
        rom[86][51] = 8'd16;
        rom[86][52] = 8'd12;
        rom[86][53] = 8'd20;
        rom[86][54] = -8'd40;
        rom[86][55] = 8'd3;
        rom[86][56] = -8'd12;
        rom[86][57] = -8'd5;
        rom[86][58] = -8'd14;
        rom[86][59] = -8'd25;
        rom[86][60] = -8'd17;
        rom[86][61] = -8'd23;
        rom[86][62] = -8'd37;
        rom[86][63] = -8'd12;
        rom[87][0] = 8'd30;
        rom[87][1] = 8'd17;
        rom[87][2] = -8'd26;
        rom[87][3] = -8'd9;
        rom[87][4] = 8'd4;
        rom[87][5] = 8'd24;
        rom[87][6] = 8'd10;
        rom[87][7] = 8'd5;
        rom[87][8] = -8'd13;
        rom[87][9] = 8'd1;
        rom[87][10] = -8'd3;
        rom[87][11] = 8'd37;
        rom[87][12] = 8'd52;
        rom[87][13] = -8'd18;
        rom[87][14] = -8'd25;
        rom[87][15] = -8'd36;
        rom[87][16] = -8'd5;
        rom[87][17] = -8'd18;
        rom[87][18] = 8'd33;
        rom[87][19] = 8'd3;
        rom[87][20] = -8'd2;
        rom[87][21] = -8'd21;
        rom[87][22] = 8'd52;
        rom[87][23] = -8'd38;
        rom[87][24] = 8'd27;
        rom[87][25] = 8'd18;
        rom[87][26] = -8'd53;
        rom[87][27] = 8'd34;
        rom[87][28] = -8'd69;
        rom[87][29] = -8'd9;
        rom[87][30] = -8'd16;
        rom[87][31] = 8'd46;
        rom[87][32] = 8'd13;
        rom[87][33] = 8'd4;
        rom[87][34] = 8'd17;
        rom[87][35] = 8'd37;
        rom[87][36] = 8'd8;
        rom[87][37] = 8'd0;
        rom[87][38] = 8'd51;
        rom[87][39] = 8'd11;
        rom[87][40] = 8'd33;
        rom[87][41] = 8'd20;
        rom[87][42] = 8'd32;
        rom[87][43] = -8'd11;
        rom[87][44] = 8'd31;
        rom[87][45] = -8'd21;
        rom[87][46] = 8'd15;
        rom[87][47] = 8'd13;
        rom[87][48] = -8'd6;
        rom[87][49] = -8'd52;
        rom[87][50] = -8'd29;
        rom[87][51] = -8'd42;
        rom[87][52] = 8'd18;
        rom[87][53] = -8'd19;
        rom[87][54] = -8'd5;
        rom[87][55] = -8'd6;
        rom[87][56] = -8'd3;
        rom[87][57] = -8'd1;
        rom[87][58] = 8'd31;
        rom[87][59] = 8'd17;
        rom[87][60] = 8'd13;
        rom[87][61] = -8'd53;
        rom[87][62] = -8'd15;
        rom[87][63] = -8'd3;
        rom[88][0] = -8'd34;
        rom[88][1] = 8'd7;
        rom[88][2] = 8'd18;
        rom[88][3] = -8'd35;
        rom[88][4] = -8'd5;
        rom[88][5] = 8'd5;
        rom[88][6] = 8'd11;
        rom[88][7] = 8'd33;
        rom[88][8] = 8'd23;
        rom[88][9] = -8'd2;
        rom[88][10] = 8'd3;
        rom[88][11] = 8'd32;
        rom[88][12] = 8'd15;
        rom[88][13] = 8'd2;
        rom[88][14] = 8'd6;
        rom[88][15] = -8'd11;
        rom[88][16] = 8'd21;
        rom[88][17] = 8'd19;
        rom[88][18] = 8'd11;
        rom[88][19] = 8'd0;
        rom[88][20] = -8'd6;
        rom[88][21] = 8'd24;
        rom[88][22] = -8'd7;
        rom[88][23] = -8'd5;
        rom[88][24] = 8'd8;
        rom[88][25] = 8'd20;
        rom[88][26] = 8'd1;
        rom[88][27] = 8'd23;
        rom[88][28] = -8'd22;
        rom[88][29] = 8'd6;
        rom[88][30] = 8'd20;
        rom[88][31] = -8'd1;
        rom[88][32] = -8'd1;
        rom[88][33] = -8'd10;
        rom[88][34] = 8'd26;
        rom[88][35] = 8'd5;
        rom[88][36] = 8'd19;
        rom[88][37] = -8'd19;
        rom[88][38] = 8'd26;
        rom[88][39] = 8'd8;
        rom[88][40] = 8'd41;
        rom[88][41] = 8'd28;
        rom[88][42] = 8'd15;
        rom[88][43] = 8'd28;
        rom[88][44] = 8'd14;
        rom[88][45] = 8'd19;
        rom[88][46] = 8'd10;
        rom[88][47] = -8'd37;
        rom[88][48] = -8'd9;
        rom[88][49] = 8'd10;
        rom[88][50] = -8'd5;
        rom[88][51] = 8'd9;
        rom[88][52] = 8'd4;
        rom[88][53] = -8'd8;
        rom[88][54] = -8'd15;
        rom[88][55] = 8'd9;
        rom[88][56] = 8'd26;
        rom[88][57] = -8'd1;
        rom[88][58] = 8'd4;
        rom[88][59] = -8'd9;
        rom[88][60] = 8'd5;
        rom[88][61] = -8'd9;
        rom[88][62] = 8'd6;
        rom[88][63] = 8'd2;
        rom[89][0] = 8'd19;
        rom[89][1] = 8'd20;
        rom[89][2] = -8'd41;
        rom[89][3] = 8'd13;
        rom[89][4] = 8'd51;
        rom[89][5] = 8'd12;
        rom[89][6] = 8'd26;
        rom[89][7] = 8'd12;
        rom[89][8] = 8'd9;
        rom[89][9] = 8'd0;
        rom[89][10] = -8'd12;
        rom[89][11] = -8'd3;
        rom[89][12] = 8'd28;
        rom[89][13] = -8'd37;
        rom[89][14] = -8'd3;
        rom[89][15] = 8'd3;
        rom[89][16] = 8'd37;
        rom[89][17] = 8'd21;
        rom[89][18] = -8'd11;
        rom[89][19] = 8'd17;
        rom[89][20] = 8'd4;
        rom[89][21] = 8'd18;
        rom[89][22] = -8'd28;
        rom[89][23] = 8'd11;
        rom[89][24] = -8'd20;
        rom[89][25] = 8'd15;
        rom[89][26] = 8'd52;
        rom[89][27] = -8'd44;
        rom[89][28] = -8'd3;
        rom[89][29] = -8'd20;
        rom[89][30] = -8'd27;
        rom[89][31] = -8'd5;
        rom[89][32] = 8'd8;
        rom[89][33] = -8'd8;
        rom[89][34] = -8'd10;
        rom[89][35] = 8'd3;
        rom[89][36] = 8'd23;
        rom[89][37] = 8'd32;
        rom[89][38] = -8'd4;
        rom[89][39] = -8'd20;
        rom[89][40] = 8'd24;
        rom[89][41] = 8'd41;
        rom[89][42] = -8'd34;
        rom[89][43] = -8'd24;
        rom[89][44] = -8'd21;
        rom[89][45] = 8'd21;
        rom[89][46] = -8'd5;
        rom[89][47] = -8'd23;
        rom[89][48] = -8'd37;
        rom[89][49] = -8'd20;
        rom[89][50] = -8'd2;
        rom[89][51] = 8'd36;
        rom[89][52] = -8'd45;
        rom[89][53] = 8'd7;
        rom[89][54] = -8'd1;
        rom[89][55] = 8'd2;
        rom[89][56] = 8'd37;
        rom[89][57] = 8'd3;
        rom[89][58] = 8'd28;
        rom[89][59] = 8'd18;
        rom[89][60] = 8'd39;
        rom[89][61] = 8'd34;
        rom[89][62] = -8'd31;
        rom[89][63] = -8'd14;
        rom[90][0] = -8'd16;
        rom[90][1] = -8'd12;
        rom[90][2] = 8'd8;
        rom[90][3] = -8'd51;
        rom[90][4] = -8'd9;
        rom[90][5] = 8'd25;
        rom[90][6] = 8'd5;
        rom[90][7] = 8'd4;
        rom[90][8] = 8'd6;
        rom[90][9] = -8'd2;
        rom[90][10] = 8'd10;
        rom[90][11] = -8'd10;
        rom[90][12] = -8'd22;
        rom[90][13] = 8'd5;
        rom[90][14] = 8'd4;
        rom[90][15] = -8'd42;
        rom[90][16] = -8'd10;
        rom[90][17] = 8'd30;
        rom[90][18] = -8'd48;
        rom[90][19] = 8'd38;
        rom[90][20] = -8'd6;
        rom[90][21] = -8'd21;
        rom[90][22] = -8'd7;
        rom[90][23] = 8'd9;
        rom[90][24] = -8'd17;
        rom[90][25] = -8'd8;
        rom[90][26] = 8'd3;
        rom[90][27] = 8'd6;
        rom[90][28] = -8'd2;
        rom[90][29] = -8'd51;
        rom[90][30] = 8'd19;
        rom[90][31] = -8'd6;
        rom[90][32] = -8'd17;
        rom[90][33] = 8'd2;
        rom[90][34] = -8'd16;
        rom[90][35] = -8'd26;
        rom[90][36] = 8'd10;
        rom[90][37] = -8'd6;
        rom[90][38] = 8'd0;
        rom[90][39] = 8'd33;
        rom[90][40] = 8'd15;
        rom[90][41] = -8'd4;
        rom[90][42] = -8'd1;
        rom[90][43] = -8'd4;
        rom[90][44] = 8'd29;
        rom[90][45] = 8'd0;
        rom[90][46] = 8'd44;
        rom[90][47] = -8'd38;
        rom[90][48] = -8'd44;
        rom[90][49] = -8'd11;
        rom[90][50] = -8'd13;
        rom[90][51] = -8'd12;
        rom[90][52] = 8'd9;
        rom[90][53] = -8'd21;
        rom[90][54] = -8'd90;
        rom[90][55] = -8'd36;
        rom[90][56] = 8'd9;
        rom[90][57] = -8'd57;
        rom[90][58] = 8'd7;
        rom[90][59] = -8'd12;
        rom[90][60] = -8'd27;
        rom[90][61] = -8'd24;
        rom[90][62] = -8'd20;
        rom[90][63] = 8'd1;
        rom[91][0] = -8'd6;
        rom[91][1] = -8'd22;
        rom[91][2] = 8'd39;
        rom[91][3] = -8'd11;
        rom[91][4] = 8'd59;
        rom[91][5] = 8'd4;
        rom[91][6] = 8'd3;
        rom[91][7] = 8'd28;
        rom[91][8] = 8'd35;
        rom[91][9] = 8'd8;
        rom[91][10] = -8'd63;
        rom[91][11] = -8'd12;
        rom[91][12] = -8'd42;
        rom[91][13] = -8'd8;
        rom[91][14] = 8'd14;
        rom[91][15] = 8'd1;
        rom[91][16] = 8'd2;
        rom[91][17] = -8'd27;
        rom[91][18] = 8'd9;
        rom[91][19] = -8'd14;
        rom[91][20] = 8'd8;
        rom[91][21] = -8'd26;
        rom[91][22] = 8'd30;
        rom[91][23] = 8'd28;
        rom[91][24] = 8'd27;
        rom[91][25] = -8'd21;
        rom[91][26] = 8'd14;
        rom[91][27] = -8'd30;
        rom[91][28] = 8'd25;
        rom[91][29] = -8'd1;
        rom[91][30] = 8'd1;
        rom[91][31] = 8'd0;
        rom[91][32] = -8'd12;
        rom[91][33] = -8'd29;
        rom[91][34] = -8'd10;
        rom[91][35] = 8'd25;
        rom[91][36] = -8'd24;
        rom[91][37] = -8'd3;
        rom[91][38] = 8'd3;
        rom[91][39] = -8'd28;
        rom[91][40] = -8'd5;
        rom[91][41] = 8'd25;
        rom[91][42] = -8'd47;
        rom[91][43] = 8'd29;
        rom[91][44] = 8'd6;
        rom[91][45] = 8'd25;
        rom[91][46] = 8'd8;
        rom[91][47] = -8'd3;
        rom[91][48] = 8'd18;
        rom[91][49] = -8'd11;
        rom[91][50] = 8'd35;
        rom[91][51] = 8'd43;
        rom[91][52] = 8'd16;
        rom[91][53] = 8'd40;
        rom[91][54] = 8'd49;
        rom[91][55] = 8'd19;
        rom[91][56] = 8'd51;
        rom[91][57] = 8'd3;
        rom[91][58] = 8'd10;
        rom[91][59] = -8'd26;
        rom[91][60] = 8'd29;
        rom[91][61] = 8'd19;
        rom[91][62] = -8'd40;
        rom[91][63] = -8'd5;
        rom[92][0] = -8'd6;
        rom[92][1] = 8'd19;
        rom[92][2] = 8'd18;
        rom[92][3] = -8'd43;
        rom[92][4] = 8'd5;
        rom[92][5] = -8'd56;
        rom[92][6] = 8'd49;
        rom[92][7] = 8'd28;
        rom[92][8] = -8'd14;
        rom[92][9] = 8'd23;
        rom[92][10] = 8'd7;
        rom[92][11] = -8'd2;
        rom[92][12] = -8'd52;
        rom[92][13] = -8'd7;
        rom[92][14] = 8'd16;
        rom[92][15] = -8'd35;
        rom[92][16] = -8'd53;
        rom[92][17] = 8'd17;
        rom[92][18] = -8'd19;
        rom[92][19] = -8'd29;
        rom[92][20] = -8'd5;
        rom[92][21] = 8'd35;
        rom[92][22] = -8'd2;
        rom[92][23] = 8'd21;
        rom[92][24] = -8'd3;
        rom[92][25] = 8'd19;
        rom[92][26] = -8'd51;
        rom[92][27] = 8'd12;
        rom[92][28] = -8'd34;
        rom[92][29] = 8'd30;
        rom[92][30] = -8'd20;
        rom[92][31] = 8'd4;
        rom[92][32] = -8'd10;
        rom[92][33] = -8'd22;
        rom[92][34] = -8'd2;
        rom[92][35] = -8'd3;
        rom[92][36] = 8'd10;
        rom[92][37] = -8'd1;
        rom[92][38] = 8'd7;
        rom[92][39] = -8'd6;
        rom[92][40] = -8'd35;
        rom[92][41] = 8'd54;
        rom[92][42] = -8'd39;
        rom[92][43] = 8'd9;
        rom[92][44] = -8'd10;
        rom[92][45] = 8'd22;
        rom[92][46] = -8'd15;
        rom[92][47] = -8'd25;
        rom[92][48] = -8'd34;
        rom[92][49] = 8'd17;
        rom[92][50] = 8'd12;
        rom[92][51] = 8'd21;
        rom[92][52] = -8'd53;
        rom[92][53] = -8'd44;
        rom[92][54] = -8'd29;
        rom[92][55] = 8'd17;
        rom[92][56] = 8'd39;
        rom[92][57] = 8'd47;
        rom[92][58] = 8'd11;
        rom[92][59] = -8'd32;
        rom[92][60] = 8'd15;
        rom[92][61] = 8'd10;
        rom[92][62] = 8'd7;
        rom[92][63] = 8'd15;
        rom[93][0] = 8'd3;
        rom[93][1] = -8'd15;
        rom[93][2] = -8'd68;
        rom[93][3] = -8'd28;
        rom[93][4] = -8'd34;
        rom[93][5] = -8'd21;
        rom[93][6] = 8'd7;
        rom[93][7] = 8'd23;
        rom[93][8] = -8'd7;
        rom[93][9] = -8'd12;
        rom[93][10] = 8'd54;
        rom[93][11] = 8'd7;
        rom[93][12] = -8'd30;
        rom[93][13] = -8'd60;
        rom[93][14] = 8'd5;
        rom[93][15] = 8'd4;
        rom[93][16] = -8'd6;
        rom[93][17] = 8'd26;
        rom[93][18] = 8'd0;
        rom[93][19] = -8'd40;
        rom[93][20] = -8'd11;
        rom[93][21] = 8'd6;
        rom[93][22] = -8'd17;
        rom[93][23] = -8'd59;
        rom[93][24] = -8'd44;
        rom[93][25] = 8'd1;
        rom[93][26] = -8'd32;
        rom[93][27] = -8'd4;
        rom[93][28] = 8'd43;
        rom[93][29] = 8'd6;
        rom[93][30] = -8'd23;
        rom[93][31] = 8'd2;
        rom[93][32] = -8'd18;
        rom[93][33] = -8'd65;
        rom[93][34] = -8'd38;
        rom[93][35] = 8'd24;
        rom[93][36] = 8'd13;
        rom[93][37] = -8'd5;
        rom[93][38] = -8'd54;
        rom[93][39] = -8'd44;
        rom[93][40] = -8'd23;
        rom[93][41] = 8'd23;
        rom[93][42] = -8'd26;
        rom[93][43] = -8'd86;
        rom[93][44] = -8'd23;
        rom[93][45] = 8'd17;
        rom[93][46] = -8'd55;
        rom[93][47] = 8'd21;
        rom[93][48] = 8'd11;
        rom[93][49] = -8'd29;
        rom[93][50] = -8'd28;
        rom[93][51] = 8'd23;
        rom[93][52] = -8'd57;
        rom[93][53] = -8'd57;
        rom[93][54] = -8'd14;
        rom[93][55] = -8'd25;
        rom[93][56] = -8'd36;
        rom[93][57] = -8'd7;
        rom[93][58] = -8'd58;
        rom[93][59] = -8'd87;
        rom[93][60] = 8'd28;
        rom[93][61] = 8'd15;
        rom[93][62] = -8'd1;
        rom[93][63] = -8'd1;
        rom[94][0] = -8'd22;
        rom[94][1] = -8'd8;
        rom[94][2] = -8'd14;
        rom[94][3] = 8'd53;
        rom[94][4] = 8'd7;
        rom[94][5] = -8'd5;
        rom[94][6] = 8'd21;
        rom[94][7] = -8'd12;
        rom[94][8] = 8'd6;
        rom[94][9] = 8'd17;
        rom[94][10] = 8'd12;
        rom[94][11] = 8'd40;
        rom[94][12] = -8'd23;
        rom[94][13] = 8'd11;
        rom[94][14] = -8'd26;
        rom[94][15] = -8'd16;
        rom[94][16] = -8'd11;
        rom[94][17] = 8'd8;
        rom[94][18] = 8'd18;
        rom[94][19] = 8'd2;
        rom[94][20] = -8'd10;
        rom[94][21] = -8'd12;
        rom[94][22] = 8'd12;
        rom[94][23] = -8'd25;
        rom[94][24] = -8'd12;
        rom[94][25] = -8'd33;
        rom[94][26] = 8'd4;
        rom[94][27] = -8'd34;
        rom[94][28] = -8'd22;
        rom[94][29] = 8'd24;
        rom[94][30] = 8'd38;
        rom[94][31] = 8'd0;
        rom[94][32] = 8'd3;
        rom[94][33] = -8'd15;
        rom[94][34] = 8'd4;
        rom[94][35] = -8'd7;
        rom[94][36] = 8'd38;
        rom[94][37] = 8'd25;
        rom[94][38] = 8'd44;
        rom[94][39] = 8'd7;
        rom[94][40] = -8'd5;
        rom[94][41] = -8'd2;
        rom[94][42] = 8'd0;
        rom[94][43] = -8'd17;
        rom[94][44] = 8'd5;
        rom[94][45] = 8'd36;
        rom[94][46] = -8'd18;
        rom[94][47] = 8'd32;
        rom[94][48] = -8'd45;
        rom[94][49] = -8'd9;
        rom[94][50] = -8'd25;
        rom[94][51] = -8'd44;
        rom[94][52] = -8'd6;
        rom[94][53] = 8'd9;
        rom[94][54] = -8'd35;
        rom[94][55] = 8'd11;
        rom[94][56] = 8'd23;
        rom[94][57] = 8'd3;
        rom[94][58] = -8'd100;
        rom[94][59] = 8'd0;
        rom[94][60] = -8'd11;
        rom[94][61] = -8'd12;
        rom[94][62] = -8'd36;
        rom[94][63] = -8'd13;
        rom[95][0] = 8'd10;
        rom[95][1] = -8'd14;
        rom[95][2] = 8'd17;
        rom[95][3] = -8'd32;
        rom[95][4] = -8'd7;
        rom[95][5] = -8'd25;
        rom[95][6] = 8'd4;
        rom[95][7] = 8'd33;
        rom[95][8] = 8'd6;
        rom[95][9] = -8'd8;
        rom[95][10] = -8'd72;
        rom[95][11] = -8'd31;
        rom[95][12] = -8'd6;
        rom[95][13] = -8'd25;
        rom[95][14] = -8'd29;
        rom[95][15] = 8'd11;
        rom[95][16] = 8'd7;
        rom[95][17] = 8'd1;
        rom[95][18] = -8'd37;
        rom[95][19] = 8'd46;
        rom[95][20] = 8'd0;
        rom[95][21] = -8'd24;
        rom[95][22] = 8'd5;
        rom[95][23] = -8'd41;
        rom[95][24] = -8'd37;
        rom[95][25] = 8'd17;
        rom[95][26] = -8'd28;
        rom[95][27] = -8'd33;
        rom[95][28] = 8'd29;
        rom[95][29] = -8'd28;
        rom[95][30] = -8'd24;
        rom[95][31] = -8'd9;
        rom[95][32] = 8'd31;
        rom[95][33] = 8'd25;
        rom[95][34] = -8'd5;
        rom[95][35] = -8'd10;
        rom[95][36] = 8'd16;
        rom[95][37] = 8'd18;
        rom[95][38] = 8'd26;
        rom[95][39] = -8'd1;
        rom[95][40] = 8'd17;
        rom[95][41] = -8'd24;
        rom[95][42] = 8'd24;
        rom[95][43] = 8'd19;
        rom[95][44] = 8'd4;
        rom[95][45] = -8'd33;
        rom[95][46] = 8'd25;
        rom[95][47] = -8'd55;
        rom[95][48] = 8'd65;
        rom[95][49] = 8'd21;
        rom[95][50] = 8'd12;
        rom[95][51] = 8'd4;
        rom[95][52] = -8'd36;
        rom[95][53] = -8'd10;
        rom[95][54] = 8'd29;
        rom[95][55] = 8'd11;
        rom[95][56] = -8'd4;
        rom[95][57] = -8'd32;
        rom[95][58] = 8'd1;
        rom[95][59] = -8'd20;
        rom[95][60] = 8'd15;
        rom[95][61] = 8'd13;
        rom[95][62] = 8'd25;
        rom[95][63] = -8'd1;
        rom[96][0] = -8'd18;
        rom[96][1] = -8'd8;
        rom[96][2] = 8'd0;
        rom[96][3] = 8'd5;
        rom[96][4] = 8'd12;
        rom[96][5] = 8'd9;
        rom[96][6] = 8'd33;
        rom[96][7] = -8'd5;
        rom[96][8] = -8'd16;
        rom[96][9] = 8'd8;
        rom[96][10] = -8'd2;
        rom[96][11] = -8'd25;
        rom[96][12] = 8'd14;
        rom[96][13] = -8'd16;
        rom[96][14] = 8'd34;
        rom[96][15] = -8'd3;
        rom[96][16] = 8'd15;
        rom[96][17] = -8'd4;
        rom[96][18] = 8'd12;
        rom[96][19] = -8'd14;
        rom[96][20] = 8'd5;
        rom[96][21] = -8'd11;
        rom[96][22] = 8'd33;
        rom[96][23] = -8'd7;
        rom[96][24] = -8'd50;
        rom[96][25] = -8'd7;
        rom[96][26] = -8'd6;
        rom[96][27] = -8'd33;
        rom[96][28] = -8'd1;
        rom[96][29] = -8'd41;
        rom[96][30] = -8'd45;
        rom[96][31] = -8'd25;
        rom[96][32] = 8'd18;
        rom[96][33] = 8'd14;
        rom[96][34] = -8'd73;
        rom[96][35] = 8'd0;
        rom[96][36] = 8'd14;
        rom[96][37] = 8'd15;
        rom[96][38] = 8'd15;
        rom[96][39] = -8'd65;
        rom[96][40] = 8'd7;
        rom[96][41] = -8'd14;
        rom[96][42] = 8'd15;
        rom[96][43] = -8'd22;
        rom[96][44] = -8'd5;
        rom[96][45] = 8'd15;
        rom[96][46] = 8'd20;
        rom[96][47] = -8'd12;
        rom[96][48] = -8'd41;
        rom[96][49] = 8'd2;
        rom[96][50] = 8'd0;
        rom[96][51] = 8'd29;
        rom[96][52] = 8'd22;
        rom[96][53] = -8'd51;
        rom[96][54] = -8'd16;
        rom[96][55] = -8'd21;
        rom[96][56] = -8'd3;
        rom[96][57] = -8'd21;
        rom[96][58] = -8'd39;
        rom[96][59] = -8'd18;
        rom[96][60] = -8'd19;
        rom[96][61] = -8'd43;
        rom[96][62] = -8'd36;
        rom[96][63] = -8'd39;
        rom[97][0] = -8'd33;
        rom[97][1] = 8'd27;
        rom[97][2] = -8'd19;
        rom[97][3] = -8'd30;
        rom[97][4] = -8'd12;
        rom[97][5] = -8'd1;
        rom[97][6] = -8'd66;
        rom[97][7] = 8'd13;
        rom[97][8] = 8'd17;
        rom[97][9] = -8'd21;
        rom[97][10] = 8'd38;
        rom[97][11] = 8'd4;
        rom[97][12] = 8'd34;
        rom[97][13] = -8'd72;
        rom[97][14] = 8'd22;
        rom[97][15] = -8'd19;
        rom[97][16] = 8'd5;
        rom[97][17] = 8'd29;
        rom[97][18] = 8'd35;
        rom[97][19] = -8'd30;
        rom[97][20] = 8'd4;
        rom[97][21] = 8'd24;
        rom[97][22] = -8'd1;
        rom[97][23] = -8'd32;
        rom[97][24] = -8'd21;
        rom[97][25] = 8'd9;
        rom[97][26] = -8'd21;
        rom[97][27] = 8'd14;
        rom[97][28] = -8'd23;
        rom[97][29] = -8'd17;
        rom[97][30] = -8'd31;
        rom[97][31] = -8'd23;
        rom[97][32] = -8'd39;
        rom[97][33] = -8'd2;
        rom[97][34] = -8'd17;
        rom[97][35] = 8'd1;
        rom[97][36] = 8'd15;
        rom[97][37] = 8'd50;
        rom[97][38] = -8'd8;
        rom[97][39] = 8'd1;
        rom[97][40] = 8'd33;
        rom[97][41] = -8'd23;
        rom[97][42] = -8'd24;
        rom[97][43] = -8'd31;
        rom[97][44] = -8'd8;
        rom[97][45] = 8'd37;
        rom[97][46] = -8'd67;
        rom[97][47] = -8'd1;
        rom[97][48] = 8'd2;
        rom[97][49] = -8'd25;
        rom[97][50] = -8'd4;
        rom[97][51] = -8'd12;
        rom[97][52] = -8'd86;
        rom[97][53] = 8'd11;
        rom[97][54] = -8'd19;
        rom[97][55] = 8'd22;
        rom[97][56] = -8'd18;
        rom[97][57] = -8'd11;
        rom[97][58] = -8'd22;
        rom[97][59] = 8'd9;
        rom[97][60] = -8'd28;
        rom[97][61] = 8'd25;
        rom[97][62] = 8'd9;
        rom[97][63] = -8'd31;
        rom[98][0] = -8'd12;
        rom[98][1] = 8'd17;
        rom[98][2] = -8'd50;
        rom[98][3] = -8'd1;
        rom[98][4] = -8'd13;
        rom[98][5] = 8'd17;
        rom[98][6] = -8'd11;
        rom[98][7] = 8'd3;
        rom[98][8] = -8'd2;
        rom[98][9] = 8'd3;
        rom[98][10] = 8'd3;
        rom[98][11] = 8'd31;
        rom[98][12] = -8'd4;
        rom[98][13] = 8'd17;
        rom[98][14] = -8'd8;
        rom[98][15] = -8'd34;
        rom[98][16] = -8'd2;
        rom[98][17] = 8'd21;
        rom[98][18] = 8'd7;
        rom[98][19] = 8'd9;
        rom[98][20] = -8'd3;
        rom[98][21] = -8'd9;
        rom[98][22] = 8'd19;
        rom[98][23] = -8'd34;
        rom[98][24] = 8'd29;
        rom[98][25] = 8'd25;
        rom[98][26] = -8'd4;
        rom[98][27] = -8'd63;
        rom[98][28] = -8'd45;
        rom[98][29] = -8'd83;
        rom[98][30] = -8'd19;
        rom[98][31] = -8'd9;
        rom[98][32] = 8'd1;
        rom[98][33] = -8'd32;
        rom[98][34] = 8'd16;
        rom[98][35] = -8'd62;
        rom[98][36] = -8'd16;
        rom[98][37] = -8'd25;
        rom[98][38] = -8'd13;
        rom[98][39] = 8'd3;
        rom[98][40] = -8'd1;
        rom[98][41] = -8'd32;
        rom[98][42] = -8'd56;
        rom[98][43] = 8'd55;
        rom[98][44] = -8'd51;
        rom[98][45] = -8'd8;
        rom[98][46] = 8'd0;
        rom[98][47] = -8'd37;
        rom[98][48] = -8'd9;
        rom[98][49] = 8'd28;
        rom[98][50] = -8'd41;
        rom[98][51] = 8'd13;
        rom[98][52] = -8'd17;
        rom[98][53] = -8'd1;
        rom[98][54] = -8'd11;
        rom[98][55] = -8'd46;
        rom[98][56] = -8'd34;
        rom[98][57] = -8'd1;
        rom[98][58] = -8'd54;
        rom[98][59] = -8'd9;
        rom[98][60] = -8'd11;
        rom[98][61] = -8'd21;
        rom[98][62] = 8'd10;
        rom[98][63] = 8'd6;
        rom[99][0] = 8'd35;
        rom[99][1] = -8'd15;
        rom[99][2] = 8'd31;
        rom[99][3] = -8'd15;
        rom[99][4] = -8'd11;
        rom[99][5] = -8'd31;
        rom[99][6] = -8'd30;
        rom[99][7] = -8'd10;
        rom[99][8] = 8'd0;
        rom[99][9] = -8'd29;
        rom[99][10] = -8'd23;
        rom[99][11] = -8'd3;
        rom[99][12] = 8'd38;
        rom[99][13] = -8'd27;
        rom[99][14] = 8'd14;
        rom[99][15] = -8'd39;
        rom[99][16] = -8'd8;
        rom[99][17] = -8'd55;
        rom[99][18] = -8'd55;
        rom[99][19] = -8'd31;
        rom[99][20] = -8'd12;
        rom[99][21] = 8'd10;
        rom[99][22] = -8'd6;
        rom[99][23] = 8'd2;
        rom[99][24] = -8'd27;
        rom[99][25] = -8'd4;
        rom[99][26] = -8'd42;
        rom[99][27] = 8'd11;
        rom[99][28] = -8'd37;
        rom[99][29] = 8'd14;
        rom[99][30] = 8'd3;
        rom[99][31] = 8'd19;
        rom[99][32] = -8'd32;
        rom[99][33] = -8'd41;
        rom[99][34] = -8'd10;
        rom[99][35] = 8'd25;
        rom[99][36] = -8'd15;
        rom[99][37] = 8'd27;
        rom[99][38] = -8'd5;
        rom[99][39] = -8'd5;
        rom[99][40] = -8'd21;
        rom[99][41] = -8'd30;
        rom[99][42] = 8'd0;
        rom[99][43] = 8'd10;
        rom[99][44] = -8'd24;
        rom[99][45] = 8'd4;
        rom[99][46] = -8'd9;
        rom[99][47] = 8'd0;
        rom[99][48] = 8'd42;
        rom[99][49] = 8'd14;
        rom[99][50] = 8'd0;
        rom[99][51] = -8'd31;
        rom[99][52] = -8'd24;
        rom[99][53] = -8'd72;
        rom[99][54] = -8'd12;
        rom[99][55] = -8'd15;
        rom[99][56] = 8'd46;
        rom[99][57] = 8'd1;
        rom[99][58] = 8'd10;
        rom[99][59] = 8'd16;
        rom[99][60] = -8'd28;
        rom[99][61] = 8'd9;
        rom[99][62] = 8'd5;
        rom[99][63] = 8'd21;
        rom[100][0] = 8'd16;
        rom[100][1] = -8'd32;
        rom[100][2] = 8'd14;
        rom[100][3] = -8'd15;
        rom[100][4] = 8'd34;
        rom[100][5] = 8'd2;
        rom[100][6] = -8'd4;
        rom[100][7] = 8'd10;
        rom[100][8] = 8'd7;
        rom[100][9] = 8'd7;
        rom[100][10] = -8'd8;
        rom[100][11] = -8'd31;
        rom[100][12] = -8'd49;
        rom[100][13] = -8'd10;
        rom[100][14] = -8'd10;
        rom[100][15] = 8'd24;
        rom[100][16] = 8'd8;
        rom[100][17] = 8'd6;
        rom[100][18] = -8'd21;
        rom[100][19] = 8'd5;
        rom[100][20] = -8'd6;
        rom[100][21] = 8'd27;
        rom[100][22] = -8'd3;
        rom[100][23] = -8'd16;
        rom[100][24] = -8'd9;
        rom[100][25] = 8'd22;
        rom[100][26] = -8'd34;
        rom[100][27] = -8'd18;
        rom[100][28] = -8'd22;
        rom[100][29] = -8'd22;
        rom[100][30] = -8'd6;
        rom[100][31] = -8'd12;
        rom[100][32] = -8'd72;
        rom[100][33] = -8'd34;
        rom[100][34] = 8'd8;
        rom[100][35] = -8'd33;
        rom[100][36] = 8'd6;
        rom[100][37] = 8'd28;
        rom[100][38] = -8'd6;
        rom[100][39] = -8'd20;
        rom[100][40] = -8'd9;
        rom[100][41] = -8'd50;
        rom[100][42] = -8'd42;
        rom[100][43] = 8'd31;
        rom[100][44] = -8'd54;
        rom[100][45] = -8'd33;
        rom[100][46] = -8'd50;
        rom[100][47] = -8'd32;
        rom[100][48] = 8'd14;
        rom[100][49] = -8'd3;
        rom[100][50] = -8'd6;
        rom[100][51] = -8'd21;
        rom[100][52] = -8'd62;
        rom[100][53] = 8'd17;
        rom[100][54] = -8'd4;
        rom[100][55] = 8'd16;
        rom[100][56] = -8'd46;
        rom[100][57] = 8'd5;
        rom[100][58] = 8'd10;
        rom[100][59] = 8'd40;
        rom[100][60] = 8'd0;
        rom[100][61] = 8'd11;
        rom[100][62] = -8'd12;
        rom[100][63] = -8'd29;
        rom[101][0] = -8'd10;
        rom[101][1] = -8'd59;
        rom[101][2] = -8'd28;
        rom[101][3] = -8'd55;
        rom[101][4] = -8'd22;
        rom[101][5] = -8'd16;
        rom[101][6] = -8'd2;
        rom[101][7] = -8'd28;
        rom[101][8] = 8'd9;
        rom[101][9] = 8'd10;
        rom[101][10] = -8'd15;
        rom[101][11] = -8'd19;
        rom[101][12] = -8'd78;
        rom[101][13] = 8'd1;
        rom[101][14] = 8'd18;
        rom[101][15] = -8'd1;
        rom[101][16] = -8'd15;
        rom[101][17] = -8'd2;
        rom[101][18] = 8'd13;
        rom[101][19] = -8'd41;
        rom[101][20] = 8'd8;
        rom[101][21] = -8'd17;
        rom[101][22] = -8'd14;
        rom[101][23] = -8'd21;
        rom[101][24] = 8'd12;
        rom[101][25] = 8'd4;
        rom[101][26] = -8'd4;
        rom[101][27] = 8'd15;
        rom[101][28] = -8'd13;
        rom[101][29] = 8'd14;
        rom[101][30] = -8'd37;
        rom[101][31] = -8'd37;
        rom[101][32] = -8'd63;
        rom[101][33] = -8'd50;
        rom[101][34] = -8'd39;
        rom[101][35] = 8'd9;
        rom[101][36] = -8'd7;
        rom[101][37] = -8'd34;
        rom[101][38] = -8'd61;
        rom[101][39] = -8'd14;
        rom[101][40] = 8'd30;
        rom[101][41] = 8'd4;
        rom[101][42] = -8'd34;
        rom[101][43] = 8'd3;
        rom[101][44] = -8'd51;
        rom[101][45] = -8'd27;
        rom[101][46] = -8'd59;
        rom[101][47] = -8'd15;
        rom[101][48] = -8'd9;
        rom[101][49] = 8'd1;
        rom[101][50] = 8'd11;
        rom[101][51] = 8'd19;
        rom[101][52] = 8'd26;
        rom[101][53] = 8'd28;
        rom[101][54] = -8'd6;
        rom[101][55] = 8'd1;
        rom[101][56] = -8'd62;
        rom[101][57] = 8'd22;
        rom[101][58] = -8'd27;
        rom[101][59] = -8'd27;
        rom[101][60] = -8'd24;
        rom[101][61] = 8'd9;
        rom[101][62] = -8'd4;
        rom[101][63] = -8'd39;
        rom[102][0] = 8'd10;
        rom[102][1] = -8'd14;
        rom[102][2] = 8'd25;
        rom[102][3] = -8'd10;
        rom[102][4] = -8'd10;
        rom[102][5] = -8'd10;
        rom[102][6] = 8'd37;
        rom[102][7] = 8'd45;
        rom[102][8] = -8'd27;
        rom[102][9] = 8'd46;
        rom[102][10] = -8'd14;
        rom[102][11] = 8'd2;
        rom[102][12] = -8'd66;
        rom[102][13] = -8'd32;
        rom[102][14] = -8'd19;
        rom[102][15] = -8'd17;
        rom[102][16] = 8'd27;
        rom[102][17] = -8'd14;
        rom[102][18] = -8'd11;
        rom[102][19] = -8'd7;
        rom[102][20] = -8'd2;
        rom[102][21] = -8'd15;
        rom[102][22] = -8'd41;
        rom[102][23] = 8'd29;
        rom[102][24] = -8'd13;
        rom[102][25] = 8'd31;
        rom[102][26] = 8'd51;
        rom[102][27] = 8'd3;
        rom[102][28] = 8'd40;
        rom[102][29] = 8'd11;
        rom[102][30] = 8'd28;
        rom[102][31] = 8'd4;
        rom[102][32] = 8'd0;
        rom[102][33] = -8'd36;
        rom[102][34] = -8'd16;
        rom[102][35] = 8'd18;
        rom[102][36] = -8'd10;
        rom[102][37] = 8'd1;
        rom[102][38] = -8'd5;
        rom[102][39] = -8'd60;
        rom[102][40] = -8'd3;
        rom[102][41] = -8'd61;
        rom[102][42] = -8'd9;
        rom[102][43] = 8'd51;
        rom[102][44] = 8'd18;
        rom[102][45] = -8'd44;
        rom[102][46] = -8'd46;
        rom[102][47] = -8'd10;
        rom[102][48] = 8'd6;
        rom[102][49] = -8'd53;
        rom[102][50] = -8'd56;
        rom[102][51] = 8'd7;
        rom[102][52] = 8'd11;
        rom[102][53] = 8'd9;
        rom[102][54] = 8'd27;
        rom[102][55] = -8'd26;
        rom[102][56] = -8'd43;
        rom[102][57] = 8'd2;
        rom[102][58] = 8'd3;
        rom[102][59] = 8'd1;
        rom[102][60] = 8'd31;
        rom[102][61] = -8'd37;
        rom[102][62] = -8'd11;
        rom[102][63] = -8'd43;
        rom[103][0] = -8'd23;
        rom[103][1] = 8'd17;
        rom[103][2] = -8'd40;
        rom[103][3] = -8'd11;
        rom[103][4] = 8'd3;
        rom[103][5] = 8'd11;
        rom[103][6] = 8'd2;
        rom[103][7] = 8'd7;
        rom[103][8] = 8'd38;
        rom[103][9] = -8'd33;
        rom[103][10] = 8'd2;
        rom[103][11] = 8'd35;
        rom[103][12] = -8'd21;
        rom[103][13] = 8'd7;
        rom[103][14] = -8'd2;
        rom[103][15] = 8'd29;
        rom[103][16] = 8'd29;
        rom[103][17] = -8'd49;
        rom[103][18] = 8'd9;
        rom[103][19] = 8'd23;
        rom[103][20] = -8'd1;
        rom[103][21] = -8'd27;
        rom[103][22] = -8'd47;
        rom[103][23] = -8'd3;
        rom[103][24] = 8'd0;
        rom[103][25] = -8'd68;
        rom[103][26] = 8'd22;
        rom[103][27] = -8'd19;
        rom[103][28] = 8'd22;
        rom[103][29] = -8'd13;
        rom[103][30] = 8'd5;
        rom[103][31] = -8'd21;
        rom[103][32] = -8'd27;
        rom[103][33] = -8'd60;
        rom[103][34] = 8'd0;
        rom[103][35] = 8'd12;
        rom[103][36] = -8'd22;
        rom[103][37] = 8'd18;
        rom[103][38] = -8'd4;
        rom[103][39] = 8'd13;
        rom[103][40] = -8'd2;
        rom[103][41] = -8'd27;
        rom[103][42] = 8'd20;
        rom[103][43] = -8'd46;
        rom[103][44] = -8'd88;
        rom[103][45] = 8'd19;
        rom[103][46] = 8'd17;
        rom[103][47] = -8'd34;
        rom[103][48] = -8'd21;
        rom[103][49] = -8'd7;
        rom[103][50] = -8'd52;
        rom[103][51] = -8'd15;
        rom[103][52] = 8'd1;
        rom[103][53] = -8'd16;
        rom[103][54] = 8'd11;
        rom[103][55] = -8'd53;
        rom[103][56] = -8'd9;
        rom[103][57] = -8'd17;
        rom[103][58] = 8'd26;
        rom[103][59] = -8'd17;
        rom[103][60] = 8'd11;
        rom[103][61] = -8'd14;
        rom[103][62] = -8'd19;
        rom[103][63] = 8'd18;
        rom[104][0] = 8'd0;
        rom[104][1] = -8'd55;
        rom[104][2] = -8'd16;
        rom[104][3] = 8'd28;
        rom[104][4] = 8'd15;
        rom[104][5] = -8'd9;
        rom[104][6] = 8'd12;
        rom[104][7] = 8'd3;
        rom[104][8] = -8'd1;
        rom[104][9] = -8'd19;
        rom[104][10] = -8'd47;
        rom[104][11] = 8'd26;
        rom[104][12] = -8'd2;
        rom[104][13] = 8'd23;
        rom[104][14] = -8'd4;
        rom[104][15] = -8'd23;
        rom[104][16] = -8'd35;
        rom[104][17] = -8'd17;
        rom[104][18] = 8'd1;
        rom[104][19] = -8'd32;
        rom[104][20] = -8'd2;
        rom[104][21] = 8'd12;
        rom[104][22] = -8'd11;
        rom[104][23] = 8'd28;
        rom[104][24] = 8'd26;
        rom[104][25] = -8'd63;
        rom[104][26] = -8'd1;
        rom[104][27] = -8'd13;
        rom[104][28] = -8'd24;
        rom[104][29] = -8'd101;
        rom[104][30] = -8'd9;
        rom[104][31] = 8'd35;
        rom[104][32] = 8'd2;
        rom[104][33] = -8'd18;
        rom[104][34] = -8'd15;
        rom[104][35] = 8'd15;
        rom[104][36] = -8'd8;
        rom[104][37] = -8'd21;
        rom[104][38] = 8'd4;
        rom[104][39] = 8'd21;
        rom[104][40] = 8'd22;
        rom[104][41] = 8'd10;
        rom[104][42] = 8'd16;
        rom[104][43] = 8'd0;
        rom[104][44] = -8'd8;
        rom[104][45] = -8'd4;
        rom[104][46] = 8'd17;
        rom[104][47] = -8'd11;
        rom[104][48] = 8'd13;
        rom[104][49] = -8'd10;
        rom[104][50] = -8'd22;
        rom[104][51] = 8'd6;
        rom[104][52] = -8'd30;
        rom[104][53] = -8'd27;
        rom[104][54] = 8'd16;
        rom[104][55] = 8'd10;
        rom[104][56] = -8'd15;
        rom[104][57] = 8'd25;
        rom[104][58] = 8'd13;
        rom[104][59] = 8'd45;
        rom[104][60] = -8'd6;
        rom[104][61] = -8'd9;
        rom[104][62] = -8'd65;
        rom[104][63] = 8'd5;
        rom[105][0] = -8'd4;
        rom[105][1] = 8'd0;
        rom[105][2] = 8'd15;
        rom[105][3] = 8'd58;
        rom[105][4] = 8'd37;
        rom[105][5] = 8'd13;
        rom[105][6] = 8'd5;
        rom[105][7] = -8'd34;
        rom[105][8] = -8'd1;
        rom[105][9] = 8'd5;
        rom[105][10] = -8'd15;
        rom[105][11] = 8'd26;
        rom[105][12] = -8'd20;
        rom[105][13] = 8'd5;
        rom[105][14] = -8'd15;
        rom[105][15] = -8'd28;
        rom[105][16] = -8'd33;
        rom[105][17] = -8'd61;
        rom[105][18] = -8'd42;
        rom[105][19] = -8'd31;
        rom[105][20] = -8'd10;
        rom[105][21] = -8'd32;
        rom[105][22] = 8'd12;
        rom[105][23] = 8'd1;
        rom[105][24] = 8'd28;
        rom[105][25] = -8'd50;
        rom[105][26] = -8'd23;
        rom[105][27] = 8'd18;
        rom[105][28] = -8'd11;
        rom[105][29] = -8'd15;
        rom[105][30] = 8'd15;
        rom[105][31] = -8'd3;
        rom[105][32] = -8'd13;
        rom[105][33] = -8'd40;
        rom[105][34] = -8'd22;
        rom[105][35] = 8'd18;
        rom[105][36] = -8'd9;
        rom[105][37] = -8'd44;
        rom[105][38] = -8'd15;
        rom[105][39] = -8'd16;
        rom[105][40] = 8'd34;
        rom[105][41] = -8'd9;
        rom[105][42] = -8'd14;
        rom[105][43] = -8'd8;
        rom[105][44] = 8'd16;
        rom[105][45] = -8'd55;
        rom[105][46] = -8'd14;
        rom[105][47] = -8'd4;
        rom[105][48] = -8'd15;
        rom[105][49] = -8'd2;
        rom[105][50] = 8'd26;
        rom[105][51] = 8'd0;
        rom[105][52] = -8'd13;
        rom[105][53] = 8'd23;
        rom[105][54] = -8'd12;
        rom[105][55] = 8'd7;
        rom[105][56] = -8'd15;
        rom[105][57] = 8'd0;
        rom[105][58] = -8'd14;
        rom[105][59] = -8'd51;
        rom[105][60] = 8'd5;
        rom[105][61] = -8'd26;
        rom[105][62] = -8'd1;
        rom[105][63] = -8'd2;
        rom[106][0] = -8'd19;
        rom[106][1] = -8'd14;
        rom[106][2] = 8'd30;
        rom[106][3] = -8'd75;
        rom[106][4] = -8'd43;
        rom[106][5] = -8'd13;
        rom[106][6] = -8'd31;
        rom[106][7] = 8'd7;
        rom[106][8] = 8'd9;
        rom[106][9] = -8'd10;
        rom[106][10] = 8'd22;
        rom[106][11] = -8'd3;
        rom[106][12] = -8'd1;
        rom[106][13] = 8'd12;
        rom[106][14] = 8'd8;
        rom[106][15] = -8'd35;
        rom[106][16] = -8'd4;
        rom[106][17] = 8'd4;
        rom[106][18] = 8'd14;
        rom[106][19] = -8'd12;
        rom[106][20] = -8'd2;
        rom[106][21] = -8'd6;
        rom[106][22] = -8'd89;
        rom[106][23] = -8'd5;
        rom[106][24] = -8'd10;
        rom[106][25] = 8'd7;
        rom[106][26] = 8'd6;
        rom[106][27] = 8'd21;
        rom[106][28] = 8'd25;
        rom[106][29] = -8'd15;
        rom[106][30] = 8'd19;
        rom[106][31] = -8'd18;
        rom[106][32] = 8'd17;
        rom[106][33] = -8'd10;
        rom[106][34] = 8'd22;
        rom[106][35] = -8'd32;
        rom[106][36] = -8'd17;
        rom[106][37] = -8'd14;
        rom[106][38] = 8'd15;
        rom[106][39] = 8'd44;
        rom[106][40] = -8'd5;
        rom[106][41] = -8'd8;
        rom[106][42] = 8'd0;
        rom[106][43] = -8'd10;
        rom[106][44] = -8'd35;
        rom[106][45] = -8'd8;
        rom[106][46] = 8'd24;
        rom[106][47] = -8'd11;
        rom[106][48] = 8'd15;
        rom[106][49] = -8'd31;
        rom[106][50] = 8'd16;
        rom[106][51] = -8'd34;
        rom[106][52] = 8'd13;
        rom[106][53] = -8'd19;
        rom[106][54] = -8'd6;
        rom[106][55] = 8'd15;
        rom[106][56] = 8'd6;
        rom[106][57] = -8'd15;
        rom[106][58] = -8'd20;
        rom[106][59] = -8'd13;
        rom[106][60] = -8'd29;
        rom[106][61] = 8'd10;
        rom[106][62] = 8'd1;
        rom[106][63] = 8'd16;
        rom[107][0] = -8'd9;
        rom[107][1] = -8'd34;
        rom[107][2] = 8'd25;
        rom[107][3] = -8'd42;
        rom[107][4] = 8'd25;
        rom[107][5] = 8'd29;
        rom[107][6] = -8'd33;
        rom[107][7] = -8'd6;
        rom[107][8] = 8'd20;
        rom[107][9] = -8'd2;
        rom[107][10] = 8'd23;
        rom[107][11] = -8'd8;
        rom[107][12] = -8'd6;
        rom[107][13] = -8'd27;
        rom[107][14] = -8'd11;
        rom[107][15] = 8'd24;
        rom[107][16] = -8'd24;
        rom[107][17] = 8'd18;
        rom[107][18] = 8'd23;
        rom[107][19] = -8'd24;
        rom[107][20] = -8'd24;
        rom[107][21] = 8'd28;
        rom[107][22] = -8'd21;
        rom[107][23] = -8'd11;
        rom[107][24] = 8'd3;
        rom[107][25] = 8'd14;
        rom[107][26] = -8'd28;
        rom[107][27] = 8'd18;
        rom[107][28] = 8'd4;
        rom[107][29] = -8'd3;
        rom[107][30] = -8'd16;
        rom[107][31] = -8'd18;
        rom[107][32] = -8'd39;
        rom[107][33] = -8'd57;
        rom[107][34] = 8'd19;
        rom[107][35] = 8'd11;
        rom[107][36] = 8'd13;
        rom[107][37] = -8'd15;
        rom[107][38] = -8'd2;
        rom[107][39] = -8'd20;
        rom[107][40] = 8'd4;
        rom[107][41] = 8'd0;
        rom[107][42] = -8'd23;
        rom[107][43] = 8'd5;
        rom[107][44] = -8'd53;
        rom[107][45] = -8'd26;
        rom[107][46] = 8'd4;
        rom[107][47] = 8'd10;
        rom[107][48] = -8'd7;
        rom[107][49] = -8'd20;
        rom[107][50] = 8'd5;
        rom[107][51] = 8'd1;
        rom[107][52] = 8'd8;
        rom[107][53] = 8'd13;
        rom[107][54] = -8'd6;
        rom[107][55] = 8'd21;
        rom[107][56] = -8'd6;
        rom[107][57] = 8'd26;
        rom[107][58] = -8'd2;
        rom[107][59] = 8'd18;
        rom[107][60] = 8'd3;
        rom[107][61] = 8'd17;
        rom[107][62] = -8'd24;
        rom[107][63] = 8'd11;
        rom[108][0] = -8'd31;
        rom[108][1] = -8'd2;
        rom[108][2] = 8'd15;
        rom[108][3] = -8'd16;
        rom[108][4] = -8'd20;
        rom[108][5] = -8'd59;
        rom[108][6] = 8'd8;
        rom[108][7] = -8'd30;
        rom[108][8] = -8'd6;
        rom[108][9] = -8'd31;
        rom[108][10] = -8'd16;
        rom[108][11] = -8'd36;
        rom[108][12] = -8'd13;
        rom[108][13] = -8'd12;
        rom[108][14] = -8'd24;
        rom[108][15] = -8'd37;
        rom[108][16] = -8'd8;
        rom[108][17] = -8'd10;
        rom[108][18] = 8'd20;
        rom[108][19] = -8'd42;
        rom[108][20] = -8'd14;
        rom[108][21] = -8'd27;
        rom[108][22] = -8'd40;
        rom[108][23] = 8'd0;
        rom[108][24] = 8'd17;
        rom[108][25] = 8'd22;
        rom[108][26] = 8'd29;
        rom[108][27] = 8'd14;
        rom[108][28] = -8'd29;
        rom[108][29] = 8'd10;
        rom[108][30] = -8'd1;
        rom[108][31] = -8'd7;
        rom[108][32] = -8'd19;
        rom[108][33] = -8'd70;
        rom[108][34] = -8'd55;
        rom[108][35] = -8'd8;
        rom[108][36] = 8'd38;
        rom[108][37] = -8'd11;
        rom[108][38] = 8'd13;
        rom[108][39] = 8'd14;
        rom[108][40] = -8'd61;
        rom[108][41] = -8'd7;
        rom[108][42] = -8'd24;
        rom[108][43] = 8'd0;
        rom[108][44] = 8'd21;
        rom[108][45] = 8'd19;
        rom[108][46] = -8'd9;
        rom[108][47] = -8'd49;
        rom[108][48] = 8'd7;
        rom[108][49] = 8'd8;
        rom[108][50] = 8'd25;
        rom[108][51] = 8'd30;
        rom[108][52] = -8'd36;
        rom[108][53] = -8'd29;
        rom[108][54] = -8'd31;
        rom[108][55] = -8'd12;
        rom[108][56] = -8'd43;
        rom[108][57] = 8'd3;
        rom[108][58] = -8'd25;
        rom[108][59] = -8'd72;
        rom[108][60] = -8'd25;
        rom[108][61] = 8'd19;
        rom[108][62] = 8'd27;
        rom[108][63] = -8'd5;
        rom[109][0] = 8'd8;
        rom[109][1] = -8'd53;
        rom[109][2] = 8'd1;
        rom[109][3] = -8'd4;
        rom[109][4] = -8'd27;
        rom[109][5] = 8'd34;
        rom[109][6] = 8'd25;
        rom[109][7] = 8'd36;
        rom[109][8] = -8'd21;
        rom[109][9] = -8'd11;
        rom[109][10] = 8'd6;
        rom[109][11] = -8'd30;
        rom[109][12] = -8'd41;
        rom[109][13] = 8'd20;
        rom[109][14] = 8'd14;
        rom[109][15] = -8'd11;
        rom[109][16] = 8'd3;
        rom[109][17] = 8'd20;
        rom[109][18] = -8'd43;
        rom[109][19] = -8'd19;
        rom[109][20] = 8'd4;
        rom[109][21] = 8'd2;
        rom[109][22] = -8'd32;
        rom[109][23] = -8'd29;
        rom[109][24] = 8'd17;
        rom[109][25] = -8'd26;
        rom[109][26] = -8'd8;
        rom[109][27] = -8'd38;
        rom[109][28] = -8'd17;
        rom[109][29] = 8'd10;
        rom[109][30] = 8'd36;
        rom[109][31] = -8'd19;
        rom[109][32] = -8'd8;
        rom[109][33] = 8'd19;
        rom[109][34] = -8'd26;
        rom[109][35] = -8'd14;
        rom[109][36] = 8'd48;
        rom[109][37] = 8'd3;
        rom[109][38] = -8'd27;
        rom[109][39] = -8'd22;
        rom[109][40] = -8'd12;
        rom[109][41] = -8'd30;
        rom[109][42] = 8'd12;
        rom[109][43] = -8'd17;
        rom[109][44] = 8'd33;
        rom[109][45] = -8'd16;
        rom[109][46] = 8'd32;
        rom[109][47] = -8'd4;
        rom[109][48] = -8'd12;
        rom[109][49] = -8'd61;
        rom[109][50] = -8'd36;
        rom[109][51] = 8'd0;
        rom[109][52] = -8'd18;
        rom[109][53] = -8'd3;
        rom[109][54] = 8'd26;
        rom[109][55] = -8'd43;
        rom[109][56] = -8'd41;
        rom[109][57] = -8'd14;
        rom[109][58] = -8'd17;
        rom[109][59] = -8'd10;
        rom[109][60] = 8'd4;
        rom[109][61] = 8'd53;
        rom[109][62] = 8'd51;
        rom[109][63] = 8'd30;
        rom[110][0] = 8'd1;
        rom[110][1] = -8'd33;
        rom[110][2] = -8'd14;
        rom[110][3] = 8'd3;
        rom[110][4] = -8'd37;
        rom[110][5] = -8'd8;
        rom[110][6] = -8'd35;
        rom[110][7] = -8'd6;
        rom[110][8] = -8'd23;
        rom[110][9] = -8'd16;
        rom[110][10] = -8'd60;
        rom[110][11] = -8'd23;
        rom[110][12] = -8'd5;
        rom[110][13] = 8'd16;
        rom[110][14] = -8'd4;
        rom[110][15] = -8'd20;
        rom[110][16] = -8'd32;
        rom[110][17] = -8'd14;
        rom[110][18] = -8'd11;
        rom[110][19] = -8'd8;
        rom[110][20] = -8'd1;
        rom[110][21] = -8'd7;
        rom[110][22] = -8'd15;
        rom[110][23] = -8'd6;
        rom[110][24] = 8'd5;
        rom[110][25] = -8'd59;
        rom[110][26] = 8'd8;
        rom[110][27] = -8'd8;
        rom[110][28] = -8'd38;
        rom[110][29] = -8'd26;
        rom[110][30] = -8'd8;
        rom[110][31] = -8'd5;
        rom[110][32] = 8'd20;
        rom[110][33] = 8'd21;
        rom[110][34] = -8'd19;
        rom[110][35] = -8'd2;
        rom[110][36] = -8'd11;
        rom[110][37] = -8'd12;
        rom[110][38] = 8'd12;
        rom[110][39] = -8'd23;
        rom[110][40] = 8'd34;
        rom[110][41] = 8'd47;
        rom[110][42] = 8'd7;
        rom[110][43] = 8'd15;
        rom[110][44] = -8'd88;
        rom[110][45] = 8'd27;
        rom[110][46] = 8'd5;
        rom[110][47] = -8'd4;
        rom[110][48] = 8'd24;
        rom[110][49] = -8'd16;
        rom[110][50] = -8'd15;
        rom[110][51] = 8'd6;
        rom[110][52] = 8'd16;
        rom[110][53] = -8'd23;
        rom[110][54] = -8'd10;
        rom[110][55] = -8'd66;
        rom[110][56] = -8'd7;
        rom[110][57] = 8'd15;
        rom[110][58] = 8'd0;
        rom[110][59] = 8'd9;
        rom[110][60] = -8'd49;
        rom[110][61] = -8'd56;
        rom[110][62] = -8'd20;
        rom[110][63] = -8'd51;
        rom[111][0] = -8'd55;
        rom[111][1] = 8'd33;
        rom[111][2] = -8'd53;
        rom[111][3] = -8'd23;
        rom[111][4] = -8'd10;
        rom[111][5] = -8'd14;
        rom[111][6] = 8'd31;
        rom[111][7] = -8'd20;
        rom[111][8] = -8'd1;
        rom[111][9] = -8'd40;
        rom[111][10] = 8'd41;
        rom[111][11] = 8'd14;
        rom[111][12] = -8'd39;
        rom[111][13] = -8'd36;
        rom[111][14] = -8'd1;
        rom[111][15] = -8'd37;
        rom[111][16] = 8'd16;
        rom[111][17] = 8'd19;
        rom[111][18] = -8'd33;
        rom[111][19] = 8'd5;
        rom[111][20] = 8'd0;
        rom[111][21] = 8'd0;
        rom[111][22] = 8'd13;
        rom[111][23] = -8'd45;
        rom[111][24] = 8'd0;
        rom[111][25] = 8'd18;
        rom[111][26] = 8'd13;
        rom[111][27] = 8'd24;
        rom[111][28] = -8'd45;
        rom[111][29] = 8'd21;
        rom[111][30] = -8'd12;
        rom[111][31] = 8'd37;
        rom[111][32] = -8'd32;
        rom[111][33] = 8'd15;
        rom[111][34] = 8'd19;
        rom[111][35] = 8'd42;
        rom[111][36] = -8'd47;
        rom[111][37] = 8'd20;
        rom[111][38] = 8'd10;
        rom[111][39] = 8'd37;
        rom[111][40] = 8'd60;
        rom[111][41] = -8'd10;
        rom[111][42] = 8'd6;
        rom[111][43] = -8'd33;
        rom[111][44] = -8'd25;
        rom[111][45] = 8'd14;
        rom[111][46] = 8'd48;
        rom[111][47] = 8'd21;
        rom[111][48] = -8'd64;
        rom[111][49] = 8'd43;
        rom[111][50] = -8'd20;
        rom[111][51] = 8'd15;
        rom[111][52] = -8'd18;
        rom[111][53] = -8'd20;
        rom[111][54] = 8'd34;
        rom[111][55] = 8'd14;
        rom[111][56] = -8'd13;
        rom[111][57] = 8'd34;
        rom[111][58] = -8'd20;
        rom[111][59] = 8'd48;
        rom[111][60] = -8'd32;
        rom[111][61] = -8'd17;
        rom[111][62] = 8'd14;
        rom[111][63] = -8'd14;
        rom[112][0] = -8'd19;
        rom[112][1] = -8'd5;
        rom[112][2] = -8'd37;
        rom[112][3] = 8'd27;
        rom[112][4] = 8'd27;
        rom[112][5] = -8'd39;
        rom[112][6] = -8'd10;
        rom[112][7] = -8'd31;
        rom[112][8] = 8'd3;
        rom[112][9] = -8'd13;
        rom[112][10] = -8'd25;
        rom[112][11] = -8'd20;
        rom[112][12] = 8'd1;
        rom[112][13] = 8'd7;
        rom[112][14] = 8'd4;
        rom[112][15] = 8'd17;
        rom[112][16] = 8'd39;
        rom[112][17] = 8'd15;
        rom[112][18] = -8'd29;
        rom[112][19] = 8'd9;
        rom[112][20] = -8'd17;
        rom[112][21] = 8'd32;
        rom[112][22] = -8'd65;
        rom[112][23] = 8'd23;
        rom[112][24] = -8'd13;
        rom[112][25] = -8'd26;
        rom[112][26] = -8'd62;
        rom[112][27] = -8'd39;
        rom[112][28] = -8'd19;
        rom[112][29] = -8'd35;
        rom[112][30] = 8'd34;
        rom[112][31] = 8'd10;
        rom[112][32] = -8'd35;
        rom[112][33] = -8'd26;
        rom[112][34] = 8'd9;
        rom[112][35] = -8'd70;
        rom[112][36] = 8'd13;
        rom[112][37] = -8'd37;
        rom[112][38] = -8'd11;
        rom[112][39] = -8'd12;
        rom[112][40] = -8'd11;
        rom[112][41] = -8'd4;
        rom[112][42] = 8'd18;
        rom[112][43] = 8'd16;
        rom[112][44] = -8'd7;
        rom[112][45] = -8'd18;
        rom[112][46] = 8'd24;
        rom[112][47] = 8'd0;
        rom[112][48] = -8'd22;
        rom[112][49] = -8'd30;
        rom[112][50] = -8'd9;
        rom[112][51] = -8'd23;
        rom[112][52] = -8'd14;
        rom[112][53] = 8'd11;
        rom[112][54] = -8'd20;
        rom[112][55] = -8'd16;
        rom[112][56] = 8'd15;
        rom[112][57] = -8'd23;
        rom[112][58] = -8'd7;
        rom[112][59] = 8'd17;
        rom[112][60] = -8'd9;
        rom[112][61] = 8'd9;
        rom[112][62] = 8'd24;
        rom[112][63] = -8'd20;
        rom[113][0] = -8'd37;
        rom[113][1] = 8'd52;
        rom[113][2] = 8'd16;
        rom[113][3] = 8'd25;
        rom[113][4] = -8'd15;
        rom[113][5] = 8'd2;
        rom[113][6] = -8'd10;
        rom[113][7] = -8'd23;
        rom[113][8] = 8'd47;
        rom[113][9] = 8'd4;
        rom[113][10] = 8'd16;
        rom[113][11] = 8'd8;
        rom[113][12] = 8'd22;
        rom[113][13] = -8'd16;
        rom[113][14] = 8'd8;
        rom[113][15] = -8'd31;
        rom[113][16] = 8'd20;
        rom[113][17] = -8'd17;
        rom[113][18] = -8'd38;
        rom[113][19] = 8'd8;
        rom[113][20] = 8'd8;
        rom[113][21] = -8'd20;
        rom[113][22] = 8'd45;
        rom[113][23] = -8'd18;
        rom[113][24] = -8'd4;
        rom[113][25] = -8'd2;
        rom[113][26] = -8'd13;
        rom[113][27] = 8'd32;
        rom[113][28] = 8'd30;
        rom[113][29] = 8'd22;
        rom[113][30] = 8'd24;
        rom[113][31] = 8'd8;
        rom[113][32] = -8'd20;
        rom[113][33] = 8'd16;
        rom[113][34] = -8'd6;
        rom[113][35] = -8'd16;
        rom[113][36] = 8'd7;
        rom[113][37] = 8'd30;
        rom[113][38] = -8'd14;
        rom[113][39] = -8'd13;
        rom[113][40] = 8'd0;
        rom[113][41] = -8'd20;
        rom[113][42] = 8'd34;
        rom[113][43] = -8'd13;
        rom[113][44] = -8'd17;
        rom[113][45] = -8'd11;
        rom[113][46] = -8'd9;
        rom[113][47] = 8'd21;
        rom[113][48] = 8'd14;
        rom[113][49] = -8'd25;
        rom[113][50] = 8'd5;
        rom[113][51] = -8'd29;
        rom[113][52] = -8'd30;
        rom[113][53] = 8'd25;
        rom[113][54] = 8'd8;
        rom[113][55] = -8'd5;
        rom[113][56] = -8'd4;
        rom[113][57] = -8'd8;
        rom[113][58] = -8'd56;
        rom[113][59] = 8'd1;
        rom[113][60] = -8'd3;
        rom[113][61] = 8'd4;
        rom[113][62] = -8'd22;
        rom[113][63] = 8'd8;
        rom[114][0] = 8'd22;
        rom[114][1] = 8'd0;
        rom[114][2] = -8'd15;
        rom[114][3] = -8'd28;
        rom[114][4] = -8'd31;
        rom[114][5] = 8'd15;
        rom[114][6] = -8'd5;
        rom[114][7] = -8'd15;
        rom[114][8] = -8'd27;
        rom[114][9] = -8'd27;
        rom[114][10] = -8'd35;
        rom[114][11] = 8'd12;
        rom[114][12] = -8'd22;
        rom[114][13] = -8'd15;
        rom[114][14] = 8'd0;
        rom[114][15] = -8'd30;
        rom[114][16] = -8'd10;
        rom[114][17] = 8'd29;
        rom[114][18] = -8'd27;
        rom[114][19] = 8'd11;
        rom[114][20] = 8'd7;
        rom[114][21] = -8'd36;
        rom[114][22] = -8'd2;
        rom[114][23] = -8'd30;
        rom[114][24] = -8'd28;
        rom[114][25] = -8'd54;
        rom[114][26] = 8'd1;
        rom[114][27] = -8'd26;
        rom[114][28] = -8'd51;
        rom[114][29] = -8'd1;
        rom[114][30] = -8'd48;
        rom[114][31] = -8'd12;
        rom[114][32] = -8'd9;
        rom[114][33] = 8'd27;
        rom[114][34] = -8'd35;
        rom[114][35] = -8'd9;
        rom[114][36] = 8'd10;
        rom[114][37] = -8'd13;
        rom[114][38] = 8'd5;
        rom[114][39] = -8'd45;
        rom[114][40] = 8'd2;
        rom[114][41] = 8'd24;
        rom[114][42] = 8'd21;
        rom[114][43] = -8'd7;
        rom[114][44] = -8'd23;
        rom[114][45] = -8'd41;
        rom[114][46] = 8'd0;
        rom[114][47] = -8'd38;
        rom[114][48] = -8'd16;
        rom[114][49] = -8'd1;
        rom[114][50] = 8'd1;
        rom[114][51] = 8'd16;
        rom[114][52] = 8'd4;
        rom[114][53] = -8'd40;
        rom[114][54] = 8'd9;
        rom[114][55] = -8'd36;
        rom[114][56] = -8'd15;
        rom[114][57] = -8'd4;
        rom[114][58] = 8'd18;
        rom[114][59] = 8'd3;
        rom[114][60] = -8'd31;
        rom[114][61] = -8'd3;
        rom[114][62] = 8'd5;
        rom[114][63] = -8'd42;
        rom[115][0] = 8'd14;
        rom[115][1] = -8'd6;
        rom[115][2] = 8'd37;
        rom[115][3] = -8'd31;
        rom[115][4] = -8'd19;
        rom[115][5] = 8'd2;
        rom[115][6] = 8'd9;
        rom[115][7] = 8'd11;
        rom[115][8] = -8'd6;
        rom[115][9] = -8'd14;
        rom[115][10] = 8'd36;
        rom[115][11] = 8'd0;
        rom[115][12] = -8'd2;
        rom[115][13] = -8'd28;
        rom[115][14] = -8'd19;
        rom[115][15] = 8'd16;
        rom[115][16] = -8'd13;
        rom[115][17] = -8'd11;
        rom[115][18] = 8'd21;
        rom[115][19] = -8'd5;
        rom[115][20] = 8'd1;
        rom[115][21] = -8'd1;
        rom[115][22] = -8'd31;
        rom[115][23] = -8'd16;
        rom[115][24] = 8'd30;
        rom[115][25] = -8'd4;
        rom[115][26] = 8'd14;
        rom[115][27] = 8'd6;
        rom[115][28] = -8'd28;
        rom[115][29] = -8'd3;
        rom[115][30] = 8'd13;
        rom[115][31] = -8'd21;
        rom[115][32] = 8'd42;
        rom[115][33] = 8'd22;
        rom[115][34] = -8'd45;
        rom[115][35] = 8'd29;
        rom[115][36] = 8'd9;
        rom[115][37] = 8'd33;
        rom[115][38] = 8'd11;
        rom[115][39] = 8'd28;
        rom[115][40] = -8'd18;
        rom[115][41] = -8'd2;
        rom[115][42] = 8'd12;
        rom[115][43] = -8'd16;
        rom[115][44] = -8'd3;
        rom[115][45] = 8'd18;
        rom[115][46] = 8'd21;
        rom[115][47] = -8'd1;
        rom[115][48] = 8'd6;
        rom[115][49] = -8'd24;
        rom[115][50] = 8'd19;
        rom[115][51] = 8'd7;
        rom[115][52] = -8'd36;
        rom[115][53] = -8'd39;
        rom[115][54] = -8'd44;
        rom[115][55] = 8'd35;
        rom[115][56] = -8'd20;
        rom[115][57] = -8'd17;
        rom[115][58] = -8'd19;
        rom[115][59] = -8'd25;
        rom[115][60] = 8'd26;
        rom[115][61] = 8'd8;
        rom[115][62] = 8'd4;
        rom[115][63] = -8'd23;
        rom[116][0] = -8'd40;
        rom[116][1] = -8'd40;
        rom[116][2] = 8'd2;
        rom[116][3] = -8'd13;
        rom[116][4] = 8'd27;
        rom[116][5] = -8'd32;
        rom[116][6] = 8'd19;
        rom[116][7] = 8'd9;
        rom[116][8] = 8'd11;
        rom[116][9] = -8'd15;
        rom[116][10] = -8'd5;
        rom[116][11] = 8'd7;
        rom[116][12] = -8'd66;
        rom[116][13] = 8'd27;
        rom[116][14] = 8'd12;
        rom[116][15] = 8'd49;
        rom[116][16] = 8'd5;
        rom[116][17] = 8'd6;
        rom[116][18] = 8'd13;
        rom[116][19] = -8'd53;
        rom[116][20] = -8'd6;
        rom[116][21] = -8'd11;
        rom[116][22] = 8'd36;
        rom[116][23] = -8'd20;
        rom[116][24] = -8'd27;
        rom[116][25] = 8'd6;
        rom[116][26] = -8'd16;
        rom[116][27] = -8'd4;
        rom[116][28] = -8'd4;
        rom[116][29] = -8'd5;
        rom[116][30] = -8'd9;
        rom[116][31] = 8'd3;
        rom[116][32] = -8'd29;
        rom[116][33] = -8'd4;
        rom[116][34] = -8'd13;
        rom[116][35] = 8'd11;
        rom[116][36] = -8'd17;
        rom[116][37] = -8'd9;
        rom[116][38] = 8'd2;
        rom[116][39] = 8'd24;
        rom[116][40] = 8'd7;
        rom[116][41] = 8'd25;
        rom[116][42] = 8'd33;
        rom[116][43] = 8'd1;
        rom[116][44] = -8'd9;
        rom[116][45] = -8'd43;
        rom[116][46] = -8'd51;
        rom[116][47] = -8'd79;
        rom[116][48] = 8'd40;
        rom[116][49] = -8'd5;
        rom[116][50] = -8'd13;
        rom[116][51] = 8'd19;
        rom[116][52] = 8'd7;
        rom[116][53] = -8'd5;
        rom[116][54] = -8'd15;
        rom[116][55] = 8'd19;
        rom[116][56] = -8'd10;
        rom[116][57] = 8'd20;
        rom[116][58] = 8'd2;
        rom[116][59] = 8'd12;
        rom[116][60] = 8'd7;
        rom[116][61] = 8'd34;
        rom[116][62] = 8'd13;
        rom[116][63] = -8'd2;
        rom[117][0] = -8'd12;
        rom[117][1] = 8'd0;
        rom[117][2] = -8'd24;
        rom[117][3] = -8'd30;
        rom[117][4] = -8'd14;
        rom[117][5] = -8'd51;
        rom[117][6] = -8'd30;
        rom[117][7] = 8'd6;
        rom[117][8] = 8'd0;
        rom[117][9] = -8'd1;
        rom[117][10] = -8'd68;
        rom[117][11] = 8'd26;
        rom[117][12] = 8'd29;
        rom[117][13] = -8'd19;
        rom[117][14] = -8'd8;
        rom[117][15] = -8'd5;
        rom[117][16] = 8'd18;
        rom[117][17] = 8'd9;
        rom[117][18] = 8'd24;
        rom[117][19] = 8'd12;
        rom[117][20] = -8'd13;
        rom[117][21] = -8'd14;
        rom[117][22] = 8'd15;
        rom[117][23] = -8'd42;
        rom[117][24] = -8'd24;
        rom[117][25] = -8'd29;
        rom[117][26] = 8'd29;
        rom[117][27] = -8'd10;
        rom[117][28] = 8'd16;
        rom[117][29] = -8'd21;
        rom[117][30] = -8'd25;
        rom[117][31] = 8'd9;
        rom[117][32] = -8'd1;
        rom[117][33] = -8'd15;
        rom[117][34] = 8'd17;
        rom[117][35] = 8'd14;
        rom[117][36] = 8'd28;
        rom[117][37] = -8'd19;
        rom[117][38] = 8'd19;
        rom[117][39] = 8'd26;
        rom[117][40] = 8'd24;
        rom[117][41] = -8'd10;
        rom[117][42] = -8'd28;
        rom[117][43] = -8'd8;
        rom[117][44] = -8'd55;
        rom[117][45] = 8'd1;
        rom[117][46] = -8'd19;
        rom[117][47] = 8'd11;
        rom[117][48] = -8'd15;
        rom[117][49] = -8'd44;
        rom[117][50] = -8'd57;
        rom[117][51] = -8'd24;
        rom[117][52] = -8'd3;
        rom[117][53] = 8'd0;
        rom[117][54] = -8'd6;
        rom[117][55] = 8'd0;
        rom[117][56] = -8'd4;
        rom[117][57] = 8'd18;
        rom[117][58] = 8'd8;
        rom[117][59] = 8'd8;
        rom[117][60] = -8'd9;
        rom[117][61] = -8'd49;
        rom[117][62] = -8'd24;
        rom[117][63] = 8'd5;
        rom[118][0] = -8'd6;
        rom[118][1] = -8'd3;
        rom[118][2] = -8'd2;
        rom[118][3] = -8'd7;
        rom[118][4] = -8'd4;
        rom[118][5] = -8'd2;
        rom[118][6] = -8'd6;
        rom[118][7] = -8'd6;
        rom[118][8] = 8'd3;
        rom[118][9] = 8'd8;
        rom[118][10] = -8'd7;
        rom[118][11] = 8'd11;
        rom[118][12] = 8'd4;
        rom[118][13] = 8'd8;
        rom[118][14] = 8'd12;
        rom[118][15] = -8'd3;
        rom[118][16] = -8'd7;
        rom[118][17] = 8'd16;
        rom[118][18] = -8'd5;
        rom[118][19] = 8'd9;
        rom[118][20] = 8'd0;
        rom[118][21] = 8'd0;
        rom[118][22] = 8'd0;
        rom[118][23] = -8'd10;
        rom[118][24] = -8'd7;
        rom[118][25] = 8'd5;
        rom[118][26] = -8'd4;
        rom[118][27] = 8'd2;
        rom[118][28] = 8'd14;
        rom[118][29] = 8'd7;
        rom[118][30] = 8'd2;
        rom[118][31] = -8'd1;
        rom[118][32] = -8'd3;
        rom[118][33] = -8'd1;
        rom[118][34] = -8'd4;
        rom[118][35] = 8'd7;
        rom[118][36] = 8'd2;
        rom[118][37] = -8'd2;
        rom[118][38] = 8'd7;
        rom[118][39] = 8'd6;
        rom[118][40] = -8'd2;
        rom[118][41] = 8'd12;
        rom[118][42] = -8'd4;
        rom[118][43] = -8'd3;
        rom[118][44] = 8'd3;
        rom[118][45] = -8'd10;
        rom[118][46] = 8'd4;
        rom[118][47] = -8'd5;
        rom[118][48] = -8'd9;
        rom[118][49] = 8'd4;
        rom[118][50] = -8'd5;
        rom[118][51] = -8'd2;
        rom[118][52] = -8'd8;
        rom[118][53] = -8'd4;
        rom[118][54] = 8'd3;
        rom[118][55] = 8'd4;
        rom[118][56] = 8'd3;
        rom[118][57] = -8'd2;
        rom[118][58] = -8'd5;
        rom[118][59] = -8'd7;
        rom[118][60] = 8'd1;
        rom[118][61] = -8'd5;
        rom[118][62] = -8'd1;
        rom[118][63] = -8'd9;
        rom[119][0] = 8'd2;
        rom[119][1] = 8'd10;
        rom[119][2] = -8'd3;
        rom[119][3] = -8'd43;
        rom[119][4] = -8'd13;
        rom[119][5] = -8'd24;
        rom[119][6] = 8'd21;
        rom[119][7] = -8'd12;
        rom[119][8] = 8'd30;
        rom[119][9] = -8'd9;
        rom[119][10] = 8'd1;
        rom[119][11] = -8'd56;
        rom[119][12] = -8'd16;
        rom[119][13] = 8'd26;
        rom[119][14] = -8'd19;
        rom[119][15] = -8'd12;
        rom[119][16] = 8'd17;
        rom[119][17] = 8'd3;
        rom[119][18] = -8'd5;
        rom[119][19] = 8'd10;
        rom[119][20] = -8'd16;
        rom[119][21] = 8'd39;
        rom[119][22] = -8'd37;
        rom[119][23] = 8'd2;
        rom[119][24] = -8'd36;
        rom[119][25] = 8'd3;
        rom[119][26] = -8'd7;
        rom[119][27] = 8'd4;
        rom[119][28] = -8'd22;
        rom[119][29] = 8'd41;
        rom[119][30] = 8'd16;
        rom[119][31] = 8'd8;
        rom[119][32] = 8'd28;
        rom[119][33] = -8'd30;
        rom[119][34] = -8'd1;
        rom[119][35] = -8'd4;
        rom[119][36] = -8'd3;
        rom[119][37] = -8'd5;
        rom[119][38] = -8'd5;
        rom[119][39] = -8'd17;
        rom[119][40] = 8'd61;
        rom[119][41] = 8'd6;
        rom[119][42] = -8'd1;
        rom[119][43] = -8'd38;
        rom[119][44] = -8'd32;
        rom[119][45] = -8'd10;
        rom[119][46] = -8'd23;
        rom[119][47] = -8'd100;
        rom[119][48] = -8'd48;
        rom[119][49] = 8'd7;
        rom[119][50] = -8'd74;
        rom[119][51] = 8'd7;
        rom[119][52] = -8'd18;
        rom[119][53] = 8'd17;
        rom[119][54] = -8'd10;
        rom[119][55] = 8'd6;
        rom[119][56] = -8'd25;
        rom[119][57] = 8'd11;
        rom[119][58] = -8'd5;
        rom[119][59] = -8'd1;
        rom[119][60] = -8'd5;
        rom[119][61] = -8'd7;
        rom[119][62] = 8'd16;
        rom[119][63] = 8'd1;
        rom[120][0] = -8'd69;
        rom[120][1] = -8'd17;
        rom[120][2] = 8'd18;
        rom[120][3] = -8'd50;
        rom[120][4] = -8'd26;
        rom[120][5] = -8'd89;
        rom[120][6] = -8'd10;
        rom[120][7] = -8'd30;
        rom[120][8] = -8'd36;
        rom[120][9] = -8'd28;
        rom[120][10] = 8'd13;
        rom[120][11] = -8'd55;
        rom[120][12] = -8'd37;
        rom[120][13] = -8'd21;
        rom[120][14] = -8'd24;
        rom[120][15] = -8'd51;
        rom[120][16] = 8'd21;
        rom[120][17] = 8'd20;
        rom[120][18] = -8'd41;
        rom[120][19] = -8'd41;
        rom[120][20] = -8'd2;
        rom[120][21] = -8'd5;
        rom[120][22] = -8'd57;
        rom[120][23] = -8'd73;
        rom[120][24] = 8'd3;
        rom[120][25] = -8'd24;
        rom[120][26] = -8'd5;
        rom[120][27] = -8'd33;
        rom[120][28] = -8'd17;
        rom[120][29] = 8'd24;
        rom[120][30] = -8'd10;
        rom[120][31] = 8'd11;
        rom[120][32] = -8'd30;
        rom[120][33] = -8'd26;
        rom[120][34] = -8'd41;
        rom[120][35] = -8'd18;
        rom[120][36] = 8'd7;
        rom[120][37] = 8'd11;
        rom[120][38] = -8'd10;
        rom[120][39] = -8'd9;
        rom[120][40] = 8'd18;
        rom[120][41] = -8'd23;
        rom[120][42] = -8'd42;
        rom[120][43] = 8'd24;
        rom[120][44] = -8'd1;
        rom[120][45] = -8'd51;
        rom[120][46] = 8'd9;
        rom[120][47] = -8'd57;
        rom[120][48] = -8'd16;
        rom[120][49] = 8'd6;
        rom[120][50] = 8'd35;
        rom[120][51] = 8'd6;
        rom[120][52] = -8'd6;
        rom[120][53] = 8'd9;
        rom[120][54] = -8'd44;
        rom[120][55] = 8'd10;
        rom[120][56] = -8'd19;
        rom[120][57] = -8'd21;
        rom[120][58] = -8'd86;
        rom[120][59] = -8'd4;
        rom[120][60] = -8'd21;
        rom[120][61] = 8'd35;
        rom[120][62] = 8'd0;
        rom[120][63] = -8'd43;
        rom[121][0] = -8'd1;
        rom[121][1] = -8'd7;
        rom[121][2] = 8'd30;
        rom[121][3] = 8'd12;
        rom[121][4] = 8'd15;
        rom[121][5] = 8'd14;
        rom[121][6] = 8'd3;
        rom[121][7] = 8'd10;
        rom[121][8] = 8'd18;
        rom[121][9] = 8'd8;
        rom[121][10] = 8'd19;
        rom[121][11] = -8'd18;
        rom[121][12] = -8'd11;
        rom[121][13] = -8'd1;
        rom[121][14] = 8'd25;
        rom[121][15] = -8'd15;
        rom[121][16] = -8'd8;
        rom[121][17] = 8'd42;
        rom[121][18] = -8'd28;
        rom[121][19] = -8'd5;
        rom[121][20] = 8'd6;
        rom[121][21] = 8'd4;
        rom[121][22] = 8'd28;
        rom[121][23] = 8'd16;
        rom[121][24] = 8'd16;
        rom[121][25] = -8'd9;
        rom[121][26] = -8'd17;
        rom[121][27] = -8'd38;
        rom[121][28] = -8'd25;
        rom[121][29] = 8'd44;
        rom[121][30] = 8'd6;
        rom[121][31] = -8'd7;
        rom[121][32] = 8'd28;
        rom[121][33] = 8'd3;
        rom[121][34] = -8'd27;
        rom[121][35] = -8'd17;
        rom[121][36] = 8'd3;
        rom[121][37] = 8'd11;
        rom[121][38] = 8'd26;
        rom[121][39] = 8'd21;
        rom[121][40] = -8'd14;
        rom[121][41] = -8'd21;
        rom[121][42] = 8'd16;
        rom[121][43] = -8'd16;
        rom[121][44] = 8'd34;
        rom[121][45] = 8'd6;
        rom[121][46] = -8'd14;
        rom[121][47] = 8'd28;
        rom[121][48] = 8'd24;
        rom[121][49] = -8'd13;
        rom[121][50] = -8'd27;
        rom[121][51] = -8'd14;
        rom[121][52] = -8'd14;
        rom[121][53] = -8'd66;
        rom[121][54] = 8'd21;
        rom[121][55] = 8'd8;
        rom[121][56] = 8'd0;
        rom[121][57] = 8'd4;
        rom[121][58] = -8'd24;
        rom[121][59] = -8'd1;
        rom[121][60] = 8'd34;
        rom[121][61] = -8'd7;
        rom[121][62] = -8'd15;
        rom[121][63] = 8'd32;
        rom[122][0] = 8'd41;
        rom[122][1] = -8'd6;
        rom[122][2] = -8'd8;
        rom[122][3] = 8'd6;
        rom[122][4] = 8'd4;
        rom[122][5] = 8'd36;
        rom[122][6] = 8'd5;
        rom[122][7] = -8'd41;
        rom[122][8] = -8'd46;
        rom[122][9] = 8'd2;
        rom[122][10] = 8'd46;
        rom[122][11] = -8'd50;
        rom[122][12] = 8'd1;
        rom[122][13] = 8'd3;
        rom[122][14] = 8'd1;
        rom[122][15] = -8'd2;
        rom[122][16] = -8'd14;
        rom[122][17] = 8'd12;
        rom[122][18] = -8'd41;
        rom[122][19] = 8'd14;
        rom[122][20] = -8'd5;
        rom[122][21] = -8'd6;
        rom[122][22] = 8'd29;
        rom[122][23] = -8'd1;
        rom[122][24] = -8'd17;
        rom[122][25] = -8'd40;
        rom[122][26] = 8'd33;
        rom[122][27] = 8'd26;
        rom[122][28] = -8'd72;
        rom[122][29] = -8'd58;
        rom[122][30] = -8'd11;
        rom[122][31] = 8'd1;
        rom[122][32] = -8'd33;
        rom[122][33] = 8'd20;
        rom[122][34] = -8'd28;
        rom[122][35] = -8'd3;
        rom[122][36] = 8'd2;
        rom[122][37] = 8'd15;
        rom[122][38] = 8'd44;
        rom[122][39] = -8'd21;
        rom[122][40] = 8'd14;
        rom[122][41] = 8'd29;
        rom[122][42] = -8'd29;
        rom[122][43] = -8'd53;
        rom[122][44] = -8'd9;
        rom[122][45] = -8'd20;
        rom[122][46] = -8'd19;
        rom[122][47] = -8'd17;
        rom[122][48] = 8'd53;
        rom[122][49] = -8'd29;
        rom[122][50] = 8'd2;
        rom[122][51] = -8'd31;
        rom[122][52] = -8'd46;
        rom[122][53] = 8'd12;
        rom[122][54] = -8'd29;
        rom[122][55] = 8'd26;
        rom[122][56] = 8'd44;
        rom[122][57] = -8'd27;
        rom[122][58] = 8'd26;
        rom[122][59] = 8'd18;
        rom[122][60] = 8'd15;
        rom[122][61] = 8'd31;
        rom[122][62] = -8'd2;
        rom[122][63] = -8'd8;
        rom[123][0] = 8'd1;
        rom[123][1] = -8'd30;
        rom[123][2] = -8'd57;
        rom[123][3] = -8'd11;
        rom[123][4] = -8'd4;
        rom[123][5] = -8'd19;
        rom[123][6] = -8'd9;
        rom[123][7] = 8'd7;
        rom[123][8] = 8'd18;
        rom[123][9] = 8'd23;
        rom[123][10] = 8'd16;
        rom[123][11] = -8'd57;
        rom[123][12] = -8'd20;
        rom[123][13] = -8'd23;
        rom[123][14] = 8'd4;
        rom[123][15] = 8'd18;
        rom[123][16] = 8'd0;
        rom[123][17] = 8'd10;
        rom[123][18] = -8'd17;
        rom[123][19] = 8'd2;
        rom[123][20] = -8'd4;
        rom[123][21] = 8'd27;
        rom[123][22] = -8'd2;
        rom[123][23] = -8'd7;
        rom[123][24] = 8'd0;
        rom[123][25] = 8'd14;
        rom[123][26] = -8'd29;
        rom[123][27] = -8'd35;
        rom[123][28] = 8'd16;
        rom[123][29] = -8'd13;
        rom[123][30] = -8'd34;
        rom[123][31] = -8'd25;
        rom[123][32] = -8'd59;
        rom[123][33] = -8'd81;
        rom[123][34] = 8'd27;
        rom[123][35] = -8'd12;
        rom[123][36] = 8'd3;
        rom[123][37] = -8'd30;
        rom[123][38] = 8'd16;
        rom[123][39] = -8'd3;
        rom[123][40] = 8'd4;
        rom[123][41] = -8'd16;
        rom[123][42] = -8'd1;
        rom[123][43] = -8'd5;
        rom[123][44] = -8'd27;
        rom[123][45] = 8'd6;
        rom[123][46] = -8'd34;
        rom[123][47] = -8'd8;
        rom[123][48] = -8'd27;
        rom[123][49] = 8'd20;
        rom[123][50] = 8'd4;
        rom[123][51] = -8'd14;
        rom[123][52] = -8'd16;
        rom[123][53] = 8'd5;
        rom[123][54] = -8'd17;
        rom[123][55] = 8'd13;
        rom[123][56] = -8'd63;
        rom[123][57] = 8'd4;
        rom[123][58] = 8'd8;
        rom[123][59] = -8'd11;
        rom[123][60] = 8'd8;
        rom[123][61] = 8'd24;
        rom[123][62] = 8'd16;
        rom[123][63] = 8'd1;
        rom[124][0] = -8'd2;
        rom[124][1] = -8'd15;
        rom[124][2] = 8'd6;
        rom[124][3] = 8'd15;
        rom[124][4] = 8'd12;
        rom[124][5] = -8'd36;
        rom[124][6] = -8'd41;
        rom[124][7] = 8'd26;
        rom[124][8] = 8'd0;
        rom[124][9] = 8'd7;
        rom[124][10] = -8'd62;
        rom[124][11] = -8'd11;
        rom[124][12] = 8'd54;
        rom[124][13] = -8'd3;
        rom[124][14] = 8'd4;
        rom[124][15] = 8'd1;
        rom[124][16] = 8'd11;
        rom[124][17] = 8'd10;
        rom[124][18] = 8'd5;
        rom[124][19] = -8'd6;
        rom[124][20] = 8'd3;
        rom[124][21] = -8'd7;
        rom[124][22] = -8'd22;
        rom[124][23] = 8'd21;
        rom[124][24] = 8'd2;
        rom[124][25] = 8'd0;
        rom[124][26] = 8'd14;
        rom[124][27] = 8'd28;
        rom[124][28] = 8'd0;
        rom[124][29] = -8'd10;
        rom[124][30] = -8'd22;
        rom[124][31] = 8'd1;
        rom[124][32] = -8'd8;
        rom[124][33] = -8'd39;
        rom[124][34] = -8'd34;
        rom[124][35] = 8'd25;
        rom[124][36] = 8'd18;
        rom[124][37] = 8'd20;
        rom[124][38] = 8'd2;
        rom[124][39] = -8'd18;
        rom[124][40] = 8'd13;
        rom[124][41] = 8'd12;
        rom[124][42] = -8'd31;
        rom[124][43] = -8'd13;
        rom[124][44] = 8'd23;
        rom[124][45] = 8'd45;
        rom[124][46] = 8'd16;
        rom[124][47] = -8'd43;
        rom[124][48] = -8'd42;
        rom[124][49] = 8'd6;
        rom[124][50] = 8'd19;
        rom[124][51] = -8'd35;
        rom[124][52] = -8'd33;
        rom[124][53] = 8'd3;
        rom[124][54] = 8'd31;
        rom[124][55] = 8'd26;
        rom[124][56] = -8'd6;
        rom[124][57] = 8'd29;
        rom[124][58] = 8'd26;
        rom[124][59] = 8'd30;
        rom[124][60] = -8'd48;
        rom[124][61] = 8'd20;
        rom[124][62] = -8'd53;
        rom[124][63] = -8'd27;
        rom[125][0] = 8'd31;
        rom[125][1] = -8'd6;
        rom[125][2] = 8'd46;
        rom[125][3] = 8'd45;
        rom[125][4] = 8'd0;
        rom[125][5] = 8'd1;
        rom[125][6] = 8'd13;
        rom[125][7] = -8'd4;
        rom[125][8] = 8'd40;
        rom[125][9] = 8'd32;
        rom[125][10] = 8'd30;
        rom[125][11] = -8'd25;
        rom[125][12] = -8'd53;
        rom[125][13] = -8'd14;
        rom[125][14] = 8'd23;
        rom[125][15] = -8'd6;
        rom[125][16] = 8'd0;
        rom[125][17] = 8'd2;
        rom[125][18] = -8'd25;
        rom[125][19] = -8'd21;
        rom[125][20] = 8'd4;
        rom[125][21] = 8'd11;
        rom[125][22] = 8'd34;
        rom[125][23] = 8'd0;
        rom[125][24] = 8'd8;
        rom[125][25] = -8'd7;
        rom[125][26] = -8'd7;
        rom[125][27] = -8'd15;
        rom[125][28] = -8'd53;
        rom[125][29] = 8'd32;
        rom[125][30] = -8'd31;
        rom[125][31] = -8'd5;
        rom[125][32] = 8'd1;
        rom[125][33] = 8'd24;
        rom[125][34] = -8'd17;
        rom[125][35] = 8'd40;
        rom[125][36] = -8'd4;
        rom[125][37] = 8'd9;
        rom[125][38] = -8'd33;
        rom[125][39] = 8'd0;
        rom[125][40] = -8'd34;
        rom[125][41] = 8'd12;
        rom[125][42] = -8'd32;
        rom[125][43] = -8'd39;
        rom[125][44] = -8'd17;
        rom[125][45] = -8'd20;
        rom[125][46] = -8'd13;
        rom[125][47] = 8'd25;
        rom[125][48] = 8'd8;
        rom[125][49] = -8'd57;
        rom[125][50] = 8'd28;
        rom[125][51] = -8'd29;
        rom[125][52] = 8'd2;
        rom[125][53] = -8'd12;
        rom[125][54] = -8'd7;
        rom[125][55] = -8'd11;
        rom[125][56] = 8'd2;
        rom[125][57] = 8'd0;
        rom[125][58] = -8'd44;
        rom[125][59] = -8'd35;
        rom[125][60] = -8'd1;
        rom[125][61] = -8'd68;
        rom[125][62] = -8'd33;
        rom[125][63] = 8'd8;
        rom[126][0] = 8'd43;
        rom[126][1] = -8'd30;
        rom[126][2] = -8'd25;
        rom[126][3] = -8'd7;
        rom[126][4] = -8'd64;
        rom[126][5] = -8'd6;
        rom[126][6] = -8'd21;
        rom[126][7] = -8'd10;
        rom[126][8] = -8'd65;
        rom[126][9] = 8'd0;
        rom[126][10] = -8'd18;
        rom[126][11] = 8'd15;
        rom[126][12] = 8'd39;
        rom[126][13] = -8'd21;
        rom[126][14] = -8'd23;
        rom[126][15] = 8'd28;
        rom[126][16] = -8'd4;
        rom[126][17] = 8'd26;
        rom[126][18] = 8'd22;
        rom[126][19] = 8'd1;
        rom[126][20] = -8'd6;
        rom[126][21] = 8'd16;
        rom[126][22] = -8'd128;
        rom[126][23] = 8'd29;
        rom[126][24] = 8'd20;
        rom[126][25] = 8'd44;
        rom[126][26] = -8'd55;
        rom[126][27] = -8'd49;
        rom[126][28] = 8'd37;
        rom[126][29] = -8'd36;
        rom[126][30] = 8'd26;
        rom[126][31] = -8'd17;
        rom[126][32] = -8'd13;
        rom[126][33] = 8'd0;
        rom[126][34] = 8'd6;
        rom[126][35] = 8'd0;
        rom[126][36] = 8'd2;
        rom[126][37] = -8'd7;
        rom[126][38] = 8'd1;
        rom[126][39] = 8'd19;
        rom[126][40] = 8'd44;
        rom[126][41] = -8'd15;
        rom[126][42] = -8'd78;
        rom[126][43] = -8'd56;
        rom[126][44] = 8'd12;
        rom[126][45] = -8'd6;
        rom[126][46] = -8'd18;
        rom[126][47] = -8'd16;
        rom[126][48] = -8'd42;
        rom[126][49] = -8'd28;
        rom[126][50] = -8'd34;
        rom[126][51] = -8'd8;
        rom[126][52] = 8'd7;
        rom[126][53] = -8'd22;
        rom[126][54] = 8'd0;
        rom[126][55] = 8'd4;
        rom[126][56] = 8'd25;
        rom[126][57] = -8'd18;
        rom[126][58] = -8'd46;
        rom[126][59] = -8'd30;
        rom[126][60] = -8'd15;
        rom[126][61] = -8'd10;
        rom[126][62] = -8'd13;
        rom[126][63] = 8'd0;
        rom[127][0] = -8'd4;
        rom[127][1] = -8'd25;
        rom[127][2] = -8'd43;
        rom[127][3] = 8'd5;
        rom[127][4] = -8'd19;
        rom[127][5] = 8'd29;
        rom[127][6] = 8'd0;
        rom[127][7] = -8'd14;
        rom[127][8] = 8'd0;
        rom[127][9] = 8'd7;
        rom[127][10] = -8'd8;
        rom[127][11] = 8'd24;
        rom[127][12] = 8'd5;
        rom[127][13] = -8'd20;
        rom[127][14] = -8'd68;
        rom[127][15] = 8'd4;
        rom[127][16] = -8'd34;
        rom[127][17] = 8'd7;
        rom[127][18] = 8'd19;
        rom[127][19] = -8'd5;
        rom[127][20] = -8'd6;
        rom[127][21] = 8'd24;
        rom[127][22] = -8'd36;
        rom[127][23] = -8'd1;
        rom[127][24] = 8'd23;
        rom[127][25] = -8'd65;
        rom[127][26] = 8'd21;
        rom[127][27] = -8'd45;
        rom[127][28] = -8'd17;
        rom[127][29] = -8'd57;
        rom[127][30] = -8'd15;
        rom[127][31] = -8'd9;
        rom[127][32] = -8'd6;
        rom[127][33] = -8'd28;
        rom[127][34] = -8'd4;
        rom[127][35] = -8'd26;
        rom[127][36] = -8'd34;
        rom[127][37] = 8'd9;
        rom[127][38] = 8'd32;
        rom[127][39] = 8'd28;
        rom[127][40] = -8'd4;
        rom[127][41] = 8'd15;
        rom[127][42] = -8'd40;
        rom[127][43] = -8'd24;
        rom[127][44] = -8'd40;
        rom[127][45] = 8'd15;
        rom[127][46] = 8'd13;
        rom[127][47] = 8'd21;
        rom[127][48] = 8'd25;
        rom[127][49] = 8'd2;
        rom[127][50] = -8'd26;
        rom[127][51] = 8'd25;
        rom[127][52] = -8'd24;
        rom[127][53] = -8'd20;
        rom[127][54] = -8'd10;
        rom[127][55] = -8'd31;
        rom[127][56] = -8'd3;
        rom[127][57] = 8'd6;
        rom[127][58] = -8'd1;
        rom[127][59] = -8'd17;
        rom[127][60] = -8'd33;
        rom[127][61] = 8'd20;
        rom[127][62] = -8'd30;
        rom[127][63] = -8'd17;
        rom[128][0] = -8'd51;
        rom[128][1] = 8'd24;
        rom[128][2] = -8'd19;
        rom[128][3] = -8'd44;
        rom[128][4] = -8'd23;
        rom[128][5] = -8'd20;
        rom[128][6] = 8'd10;
        rom[128][7] = 8'd36;
        rom[128][8] = 8'd35;
        rom[128][9] = -8'd12;
        rom[128][10] = -8'd22;
        rom[128][11] = -8'd31;
        rom[128][12] = 8'd13;
        rom[128][13] = -8'd9;
        rom[128][14] = -8'd20;
        rom[128][15] = -8'd18;
        rom[128][16] = -8'd7;
        rom[128][17] = -8'd23;
        rom[128][18] = 8'd12;
        rom[128][19] = -8'd24;
        rom[128][20] = 8'd1;
        rom[128][21] = -8'd20;
        rom[128][22] = 8'd56;
        rom[128][23] = -8'd38;
        rom[128][24] = -8'd26;
        rom[128][25] = -8'd22;
        rom[128][26] = -8'd39;
        rom[128][27] = -8'd19;
        rom[128][28] = -8'd1;
        rom[128][29] = -8'd5;
        rom[128][30] = -8'd60;
        rom[128][31] = 8'd11;
        rom[128][32] = -8'd8;
        rom[128][33] = -8'd18;
        rom[128][34] = 8'd16;
        rom[128][35] = 8'd5;
        rom[128][36] = -8'd2;
        rom[128][37] = -8'd10;
        rom[128][38] = 8'd1;
        rom[128][39] = 8'd18;
        rom[128][40] = -8'd14;
        rom[128][41] = 8'd7;
        rom[128][42] = -8'd63;
        rom[128][43] = 8'd6;
        rom[128][44] = 8'd14;
        rom[128][45] = 8'd0;
        rom[128][46] = -8'd28;
        rom[128][47] = 8'd24;
        rom[128][48] = -8'd53;
        rom[128][49] = 8'd13;
        rom[128][50] = -8'd21;
        rom[128][51] = 8'd3;
        rom[128][52] = -8'd24;
        rom[128][53] = 8'd41;
        rom[128][54] = -8'd75;
        rom[128][55] = -8'd2;
        rom[128][56] = 8'd11;
        rom[128][57] = 8'd26;
        rom[128][58] = -8'd7;
        rom[128][59] = -8'd66;
        rom[128][60] = -8'd41;
        rom[128][61] = 8'd44;
        rom[128][62] = -8'd11;
        rom[128][63] = 8'd3;
        rom[129][0] = 8'd4;
        rom[129][1] = 8'd43;
        rom[129][2] = 8'd6;
        rom[129][3] = -8'd55;
        rom[129][4] = -8'd33;
        rom[129][5] = -8'd37;
        rom[129][6] = 8'd0;
        rom[129][7] = -8'd39;
        rom[129][8] = 8'd33;
        rom[129][9] = -8'd38;
        rom[129][10] = -8'd30;
        rom[129][11] = 8'd27;
        rom[129][12] = 8'd6;
        rom[129][13] = -8'd31;
        rom[129][14] = 8'd14;
        rom[129][15] = -8'd1;
        rom[129][16] = -8'd5;
        rom[129][17] = -8'd30;
        rom[129][18] = -8'd30;
        rom[129][19] = -8'd27;
        rom[129][20] = 8'd10;
        rom[129][21] = -8'd29;
        rom[129][22] = -8'd120;
        rom[129][23] = -8'd23;
        rom[129][24] = 8'd2;
        rom[129][25] = -8'd20;
        rom[129][26] = 8'd8;
        rom[129][27] = -8'd63;
        rom[129][28] = -8'd56;
        rom[129][29] = -8'd7;
        rom[129][30] = -8'd6;
        rom[129][31] = 8'd6;
        rom[129][32] = -8'd67;
        rom[129][33] = 8'd34;
        rom[129][34] = -8'd84;
        rom[129][35] = -8'd60;
        rom[129][36] = -8'd4;
        rom[129][37] = -8'd22;
        rom[129][38] = -8'd5;
        rom[129][39] = 8'd20;
        rom[129][40] = -8'd11;
        rom[129][41] = 8'd10;
        rom[129][42] = -8'd50;
        rom[129][43] = -8'd17;
        rom[129][44] = -8'd39;
        rom[129][45] = 8'd18;
        rom[129][46] = 8'd2;
        rom[129][47] = -8'd5;
        rom[129][48] = -8'd28;
        rom[129][49] = 8'd7;
        rom[129][50] = 8'd13;
        rom[129][51] = -8'd14;
        rom[129][52] = 8'd7;
        rom[129][53] = -8'd42;
        rom[129][54] = -8'd12;
        rom[129][55] = -8'd30;
        rom[129][56] = 8'd40;
        rom[129][57] = 8'd19;
        rom[129][58] = -8'd22;
        rom[129][59] = -8'd7;
        rom[129][60] = -8'd21;
        rom[129][61] = -8'd28;
        rom[129][62] = 8'd54;
        rom[129][63] = 8'd1;
        rom[130][0] = -8'd9;
        rom[130][1] = -8'd36;
        rom[130][2] = -8'd6;
        rom[130][3] = 8'd18;
        rom[130][4] = -8'd5;
        rom[130][5] = -8'd53;
        rom[130][6] = -8'd27;
        rom[130][7] = -8'd5;
        rom[130][8] = 8'd38;
        rom[130][9] = 8'd35;
        rom[130][10] = 8'd3;
        rom[130][11] = 8'd14;
        rom[130][12] = -8'd89;
        rom[130][13] = -8'd50;
        rom[130][14] = 8'd35;
        rom[130][15] = -8'd9;
        rom[130][16] = -8'd29;
        rom[130][17] = -8'd1;
        rom[130][18] = -8'd24;
        rom[130][19] = -8'd7;
        rom[130][20] = -8'd10;
        rom[130][21] = 8'd10;
        rom[130][22] = 8'd4;
        rom[130][23] = -8'd65;
        rom[130][24] = 8'd1;
        rom[130][25] = -8'd61;
        rom[130][26] = -8'd31;
        rom[130][27] = -8'd30;
        rom[130][28] = 8'd0;
        rom[130][29] = 8'd20;
        rom[130][30] = 8'd36;
        rom[130][31] = 8'd14;
        rom[130][32] = -8'd34;
        rom[130][33] = -8'd22;
        rom[130][34] = 8'd9;
        rom[130][35] = -8'd54;
        rom[130][36] = 8'd17;
        rom[130][37] = 8'd8;
        rom[130][38] = 8'd3;
        rom[130][39] = 8'd25;
        rom[130][40] = 8'd27;
        rom[130][41] = -8'd8;
        rom[130][42] = -8'd4;
        rom[130][43] = -8'd33;
        rom[130][44] = -8'd54;
        rom[130][45] = -8'd41;
        rom[130][46] = -8'd26;
        rom[130][47] = -8'd15;
        rom[130][48] = -8'd14;
        rom[130][49] = -8'd21;
        rom[130][50] = 8'd1;
        rom[130][51] = -8'd26;
        rom[130][52] = 8'd23;
        rom[130][53] = 8'd16;
        rom[130][54] = 8'd0;
        rom[130][55] = -8'd5;
        rom[130][56] = -8'd29;
        rom[130][57] = 8'd8;
        rom[130][58] = 8'd14;
        rom[130][59] = -8'd6;
        rom[130][60] = -8'd52;
        rom[130][61] = 8'd22;
        rom[130][62] = -8'd5;
        rom[130][63] = -8'd14;
        rom[131][0] = -8'd7;
        rom[131][1] = -8'd22;
        rom[131][2] = 8'd4;
        rom[131][3] = -8'd27;
        rom[131][4] = -8'd16;
        rom[131][5] = -8'd6;
        rom[131][6] = 8'd46;
        rom[131][7] = -8'd4;
        rom[131][8] = -8'd15;
        rom[131][9] = -8'd55;
        rom[131][10] = -8'd56;
        rom[131][11] = -8'd43;
        rom[131][12] = 8'd45;
        rom[131][13] = 8'd13;
        rom[131][14] = -8'd27;
        rom[131][15] = 8'd11;
        rom[131][16] = -8'd9;
        rom[131][17] = -8'd32;
        rom[131][18] = 8'd25;
        rom[131][19] = 8'd59;
        rom[131][20] = -8'd1;
        rom[131][21] = -8'd5;
        rom[131][22] = 8'd28;
        rom[131][23] = 8'd11;
        rom[131][24] = -8'd33;
        rom[131][25] = -8'd38;
        rom[131][26] = -8'd55;
        rom[131][27] = 8'd6;
        rom[131][28] = 8'd9;
        rom[131][29] = 8'd16;
        rom[131][30] = -8'd19;
        rom[131][31] = -8'd45;
        rom[131][32] = 8'd7;
        rom[131][33] = 8'd6;
        rom[131][34] = -8'd33;
        rom[131][35] = 8'd42;
        rom[131][36] = -8'd2;
        rom[131][37] = -8'd21;
        rom[131][38] = 8'd51;
        rom[131][39] = 8'd47;
        rom[131][40] = -8'd12;
        rom[131][41] = 8'd23;
        rom[131][42] = -8'd47;
        rom[131][43] = -8'd8;
        rom[131][44] = 8'd49;
        rom[131][45] = -8'd4;
        rom[131][46] = 8'd4;
        rom[131][47] = 8'd46;
        rom[131][48] = -8'd9;
        rom[131][49] = 8'd18;
        rom[131][50] = 8'd12;
        rom[131][51] = -8'd8;
        rom[131][52] = -8'd3;
        rom[131][53] = 8'd10;
        rom[131][54] = -8'd45;
        rom[131][55] = -8'd11;
        rom[131][56] = 8'd38;
        rom[131][57] = -8'd41;
        rom[131][58] = -8'd10;
        rom[131][59] = -8'd9;
        rom[131][60] = -8'd24;
        rom[131][61] = 8'd7;
        rom[131][62] = 8'd15;
        rom[131][63] = 8'd31;
        rom[132][0] = -8'd20;
        rom[132][1] = -8'd5;
        rom[132][2] = 8'd11;
        rom[132][3] = 8'd14;
        rom[132][4] = 8'd6;
        rom[132][5] = 8'd8;
        rom[132][6] = -8'd37;
        rom[132][7] = -8'd36;
        rom[132][8] = 8'd28;
        rom[132][9] = 8'd11;
        rom[132][10] = -8'd15;
        rom[132][11] = -8'd7;
        rom[132][12] = 8'd39;
        rom[132][13] = -8'd13;
        rom[132][14] = 8'd17;
        rom[132][15] = -8'd13;
        rom[132][16] = -8'd44;
        rom[132][17] = 8'd26;
        rom[132][18] = -8'd93;
        rom[132][19] = 8'd19;
        rom[132][20] = 8'd1;
        rom[132][21] = -8'd41;
        rom[132][22] = 8'd28;
        rom[132][23] = -8'd11;
        rom[132][24] = -8'd12;
        rom[132][25] = -8'd15;
        rom[132][26] = 8'd16;
        rom[132][27] = 8'd6;
        rom[132][28] = -8'd8;
        rom[132][29] = -8'd2;
        rom[132][30] = -8'd69;
        rom[132][31] = 8'd12;
        rom[132][32] = -8'd20;
        rom[132][33] = -8'd27;
        rom[132][34] = 8'd1;
        rom[132][35] = 8'd18;
        rom[132][36] = -8'd34;
        rom[132][37] = 8'd3;
        rom[132][38] = -8'd51;
        rom[132][39] = 8'd12;
        rom[132][40] = 8'd19;
        rom[132][41] = 8'd10;
        rom[132][42] = 8'd10;
        rom[132][43] = 8'd8;
        rom[132][44] = -8'd3;
        rom[132][45] = -8'd49;
        rom[132][46] = -8'd13;
        rom[132][47] = -8'd37;
        rom[132][48] = 8'd2;
        rom[132][49] = 8'd3;
        rom[132][50] = 8'd9;
        rom[132][51] = -8'd6;
        rom[132][52] = -8'd33;
        rom[132][53] = 8'd24;
        rom[132][54] = -8'd21;
        rom[132][55] = 8'd18;
        rom[132][56] = -8'd31;
        rom[132][57] = -8'd20;
        rom[132][58] = -8'd9;
        rom[132][59] = -8'd19;
        rom[132][60] = -8'd33;
        rom[132][61] = 8'd7;
        rom[132][62] = -8'd46;
        rom[132][63] = -8'd2;
        rom[133][0] = -8'd6;
        rom[133][1] = 8'd4;
        rom[133][2] = 8'd6;
        rom[133][3] = -8'd4;
        rom[133][4] = 8'd4;
        rom[133][5] = 8'd1;
        rom[133][6] = 8'd4;
        rom[133][7] = -8'd6;
        rom[133][8] = 8'd4;
        rom[133][9] = 8'd4;
        rom[133][10] = 8'd7;
        rom[133][11] = 8'd2;
        rom[133][12] = 8'd2;
        rom[133][13] = 8'd9;
        rom[133][14] = -8'd5;
        rom[133][15] = 8'd2;
        rom[133][16] = 8'd1;
        rom[133][17] = 8'd0;
        rom[133][18] = -8'd8;
        rom[133][19] = 8'd5;
        rom[133][20] = -8'd8;
        rom[133][21] = 8'd2;
        rom[133][22] = -8'd3;
        rom[133][23] = 8'd5;
        rom[133][24] = -8'd5;
        rom[133][25] = 8'd4;
        rom[133][26] = -8'd2;
        rom[133][27] = 8'd6;
        rom[133][28] = 8'd0;
        rom[133][29] = 8'd3;
        rom[133][30] = -8'd7;
        rom[133][31] = 8'd6;
        rom[133][32] = -8'd9;
        rom[133][33] = -8'd2;
        rom[133][34] = 8'd2;
        rom[133][35] = -8'd10;
        rom[133][36] = -8'd6;
        rom[133][37] = 8'd3;
        rom[133][38] = 8'd4;
        rom[133][39] = 8'd3;
        rom[133][40] = -8'd3;
        rom[133][41] = -8'd1;
        rom[133][42] = -8'd4;
        rom[133][43] = 8'd2;
        rom[133][44] = 8'd5;
        rom[133][45] = -8'd4;
        rom[133][46] = 8'd3;
        rom[133][47] = 8'd1;
        rom[133][48] = 8'd6;
        rom[133][49] = -8'd5;
        rom[133][50] = 8'd3;
        rom[133][51] = -8'd11;
        rom[133][52] = 8'd5;
        rom[133][53] = -8'd8;
        rom[133][54] = 8'd2;
        rom[133][55] = -8'd9;
        rom[133][56] = -8'd6;
        rom[133][57] = -8'd6;
        rom[133][58] = 8'd2;
        rom[133][59] = 8'd5;
        rom[133][60] = 8'd2;
        rom[133][61] = 8'd8;
        rom[133][62] = -8'd1;
        rom[133][63] = 8'd1;
        rom[134][0] = -8'd2;
        rom[134][1] = -8'd10;
        rom[134][2] = 8'd20;
        rom[134][3] = 8'd11;
        rom[134][4] = -8'd10;
        rom[134][5] = -8'd19;
        rom[134][6] = -8'd8;
        rom[134][7] = -8'd18;
        rom[134][8] = 8'd6;
        rom[134][9] = 8'd5;
        rom[134][10] = -8'd53;
        rom[134][11] = -8'd13;
        rom[134][12] = -8'd23;
        rom[134][13] = -8'd15;
        rom[134][14] = 8'd34;
        rom[134][15] = 8'd14;
        rom[134][16] = 8'd24;
        rom[134][17] = -8'd26;
        rom[134][18] = -8'd2;
        rom[134][19] = 8'd11;
        rom[134][20] = -8'd6;
        rom[134][21] = 8'd9;
        rom[134][22] = -8'd4;
        rom[134][23] = 8'd6;
        rom[134][24] = -8'd12;
        rom[134][25] = -8'd19;
        rom[134][26] = -8'd13;
        rom[134][27] = -8'd29;
        rom[134][28] = -8'd8;
        rom[134][29] = -8'd2;
        rom[134][30] = -8'd18;
        rom[134][31] = -8'd8;
        rom[134][32] = 8'd44;
        rom[134][33] = 8'd17;
        rom[134][34] = 8'd1;
        rom[134][35] = 8'd9;
        rom[134][36] = -8'd11;
        rom[134][37] = -8'd17;
        rom[134][38] = -8'd8;
        rom[134][39] = -8'd26;
        rom[134][40] = -8'd5;
        rom[134][41] = -8'd7;
        rom[134][42] = 8'd10;
        rom[134][43] = -8'd48;
        rom[134][44] = 8'd30;
        rom[134][45] = 8'd9;
        rom[134][46] = -8'd44;
        rom[134][47] = 8'd10;
        rom[134][48] = 8'd7;
        rom[134][49] = -8'd4;
        rom[134][50] = 8'd19;
        rom[134][51] = -8'd8;
        rom[134][52] = -8'd52;
        rom[134][53] = -8'd5;
        rom[134][54] = 8'd39;
        rom[134][55] = -8'd26;
        rom[134][56] = 8'd17;
        rom[134][57] = 8'd4;
        rom[134][58] = -8'd28;
        rom[134][59] = -8'd84;
        rom[134][60] = 8'd25;
        rom[134][61] = 8'd4;
        rom[134][62] = -8'd48;
        rom[134][63] = -8'd28;
        rom[135][0] = 8'd0;
        rom[135][1] = 8'd19;
        rom[135][2] = -8'd14;
        rom[135][3] = 8'd8;
        rom[135][4] = 8'd2;
        rom[135][5] = 8'd11;
        rom[135][6] = -8'd52;
        rom[135][7] = -8'd28;
        rom[135][8] = -8'd14;
        rom[135][9] = -8'd40;
        rom[135][10] = -8'd34;
        rom[135][11] = 8'd29;
        rom[135][12] = 8'd4;
        rom[135][13] = 8'd21;
        rom[135][14] = -8'd12;
        rom[135][15] = -8'd1;
        rom[135][16] = 8'd12;
        rom[135][17] = 8'd27;
        rom[135][18] = -8'd17;
        rom[135][19] = -8'd51;
        rom[135][20] = 8'd11;
        rom[135][21] = 8'd30;
        rom[135][22] = 8'd61;
        rom[135][23] = 8'd7;
        rom[135][24] = 8'd59;
        rom[135][25] = -8'd55;
        rom[135][26] = 8'd29;
        rom[135][27] = 8'd0;
        rom[135][28] = -8'd1;
        rom[135][29] = -8'd27;
        rom[135][30] = 8'd16;
        rom[135][31] = 8'd18;
        rom[135][32] = -8'd12;
        rom[135][33] = 8'd8;
        rom[135][34] = -8'd34;
        rom[135][35] = -8'd9;
        rom[135][36] = -8'd26;
        rom[135][37] = 8'd14;
        rom[135][38] = 8'd9;
        rom[135][39] = -8'd52;
        rom[135][40] = -8'd12;
        rom[135][41] = 8'd7;
        rom[135][42] = 8'd34;
        rom[135][43] = 8'd23;
        rom[135][44] = 8'd0;
        rom[135][45] = 8'd8;
        rom[135][46] = 8'd3;
        rom[135][47] = -8'd8;
        rom[135][48] = -8'd32;
        rom[135][49] = -8'd17;
        rom[135][50] = 8'd3;
        rom[135][51] = -8'd41;
        rom[135][52] = 8'd2;
        rom[135][53] = -8'd41;
        rom[135][54] = -8'd9;
        rom[135][55] = 8'd13;
        rom[135][56] = -8'd7;
        rom[135][57] = -8'd13;
        rom[135][58] = -8'd21;
        rom[135][59] = 8'd6;
        rom[135][60] = -8'd37;
        rom[135][61] = -8'd19;
        rom[135][62] = 8'd45;
        rom[135][63] = -8'd36;
        rom[136][0] = 8'd52;
        rom[136][1] = 8'd36;
        rom[136][2] = -8'd12;
        rom[136][3] = 8'd60;
        rom[136][4] = 8'd15;
        rom[136][5] = 8'd14;
        rom[136][6] = -8'd23;
        rom[136][7] = 8'd19;
        rom[136][8] = -8'd6;
        rom[136][9] = 8'd20;
        rom[136][10] = -8'd41;
        rom[136][11] = -8'd13;
        rom[136][12] = -8'd5;
        rom[136][13] = -8'd12;
        rom[136][14] = 8'd25;
        rom[136][15] = 8'd44;
        rom[136][16] = 8'd9;
        rom[136][17] = 8'd23;
        rom[136][18] = -8'd36;
        rom[136][19] = 8'd41;
        rom[136][20] = -8'd4;
        rom[136][21] = 8'd7;
        rom[136][22] = 8'd19;
        rom[136][23] = 8'd1;
        rom[136][24] = 8'd4;
        rom[136][25] = 8'd30;
        rom[136][26] = 8'd32;
        rom[136][27] = -8'd3;
        rom[136][28] = 8'd12;
        rom[136][29] = 8'd0;
        rom[136][30] = -8'd6;
        rom[136][31] = 8'd29;
        rom[136][32] = -8'd10;
        rom[136][33] = -8'd9;
        rom[136][34] = -8'd17;
        rom[136][35] = 8'd23;
        rom[136][36] = -8'd10;
        rom[136][37] = 8'd32;
        rom[136][38] = -8'd29;
        rom[136][39] = -8'd8;
        rom[136][40] = 8'd2;
        rom[136][41] = 8'd27;
        rom[136][42] = -8'd5;
        rom[136][43] = 8'd11;
        rom[136][44] = -8'd21;
        rom[136][45] = 8'd14;
        rom[136][46] = 8'd5;
        rom[136][47] = -8'd29;
        rom[136][48] = 8'd11;
        rom[136][49] = -8'd27;
        rom[136][50] = 8'd16;
        rom[136][51] = 8'd5;
        rom[136][52] = -8'd20;
        rom[136][53] = -8'd45;
        rom[136][54] = -8'd19;
        rom[136][55] = -8'd12;
        rom[136][56] = -8'd3;
        rom[136][57] = 8'd4;
        rom[136][58] = -8'd37;
        rom[136][59] = 8'd8;
        rom[136][60] = -8'd11;
        rom[136][61] = -8'd39;
        rom[136][62] = -8'd3;
        rom[136][63] = -8'd15;
        rom[137][0] = -8'd13;
        rom[137][1] = -8'd7;
        rom[137][2] = 8'd15;
        rom[137][3] = 8'd10;
        rom[137][4] = -8'd20;
        rom[137][5] = 8'd19;
        rom[137][6] = -8'd26;
        rom[137][7] = -8'd27;
        rom[137][8] = 8'd11;
        rom[137][9] = -8'd38;
        rom[137][10] = 8'd7;
        rom[137][11] = 8'd26;
        rom[137][12] = 8'd41;
        rom[137][13] = 8'd11;
        rom[137][14] = 8'd4;
        rom[137][15] = 8'd8;
        rom[137][16] = 8'd29;
        rom[137][17] = 8'd14;
        rom[137][18] = 8'd52;
        rom[137][19] = 8'd29;
        rom[137][20] = -8'd1;
        rom[137][21] = -8'd2;
        rom[137][22] = -8'd38;
        rom[137][23] = 8'd1;
        rom[137][24] = 8'd24;
        rom[137][25] = -8'd27;
        rom[137][26] = 8'd26;
        rom[137][27] = -8'd21;
        rom[137][28] = 8'd19;
        rom[137][29] = 8'd25;
        rom[137][30] = -8'd7;
        rom[137][31] = 8'd14;
        rom[137][32] = 8'd22;
        rom[137][33] = 8'd17;
        rom[137][34] = 8'd24;
        rom[137][35] = 8'd7;
        rom[137][36] = -8'd14;
        rom[137][37] = 8'd1;
        rom[137][38] = 8'd24;
        rom[137][39] = -8'd13;
        rom[137][40] = -8'd2;
        rom[137][41] = -8'd16;
        rom[137][42] = 8'd28;
        rom[137][43] = 8'd7;
        rom[137][44] = -8'd49;
        rom[137][45] = 8'd13;
        rom[137][46] = -8'd33;
        rom[137][47] = 8'd14;
        rom[137][48] = -8'd16;
        rom[137][49] = -8'd18;
        rom[137][50] = -8'd38;
        rom[137][51] = -8'd27;
        rom[137][52] = -8'd14;
        rom[137][53] = 8'd12;
        rom[137][54] = 8'd29;
        rom[137][55] = -8'd16;
        rom[137][56] = -8'd18;
        rom[137][57] = -8'd34;
        rom[137][58] = 8'd22;
        rom[137][59] = 8'd6;
        rom[137][60] = -8'd6;
        rom[137][61] = 8'd1;
        rom[137][62] = -8'd40;
        rom[137][63] = -8'd41;
        rom[138][0] = -8'd20;
        rom[138][1] = -8'd40;
        rom[138][2] = 8'd21;
        rom[138][3] = -8'd30;
        rom[138][4] = 8'd0;
        rom[138][5] = 8'd4;
        rom[138][6] = 8'd17;
        rom[138][7] = -8'd8;
        rom[138][8] = -8'd1;
        rom[138][9] = 8'd7;
        rom[138][10] = -8'd48;
        rom[138][11] = -8'd60;
        rom[138][12] = -8'd3;
        rom[138][13] = -8'd41;
        rom[138][14] = 8'd13;
        rom[138][15] = 8'd15;
        rom[138][16] = -8'd22;
        rom[138][17] = -8'd14;
        rom[138][18] = -8'd2;
        rom[138][19] = 8'd4;
        rom[138][20] = 8'd0;
        rom[138][21] = 8'd13;
        rom[138][22] = -8'd40;
        rom[138][23] = -8'd29;
        rom[138][24] = 8'd12;
        rom[138][25] = 8'd47;
        rom[138][26] = -8'd38;
        rom[138][27] = -8'd56;
        rom[138][28] = 8'd21;
        rom[138][29] = -8'd14;
        rom[138][30] = -8'd16;
        rom[138][31] = -8'd42;
        rom[138][32] = -8'd13;
        rom[138][33] = 8'd13;
        rom[138][34] = 8'd14;
        rom[138][35] = 8'd16;
        rom[138][36] = 8'd22;
        rom[138][37] = -8'd34;
        rom[138][38] = -8'd34;
        rom[138][39] = 8'd18;
        rom[138][40] = -8'd23;
        rom[138][41] = 8'd17;
        rom[138][42] = -8'd27;
        rom[138][43] = -8'd36;
        rom[138][44] = -8'd3;
        rom[138][45] = -8'd2;
        rom[138][46] = 8'd22;
        rom[138][47] = -8'd13;
        rom[138][48] = -8'd38;
        rom[138][49] = -8'd27;
        rom[138][50] = 8'd11;
        rom[138][51] = -8'd9;
        rom[138][52] = 8'd23;
        rom[138][53] = -8'd9;
        rom[138][54] = 8'd39;
        rom[138][55] = -8'd8;
        rom[138][56] = -8'd62;
        rom[138][57] = 8'd5;
        rom[138][58] = -8'd12;
        rom[138][59] = -8'd70;
        rom[138][60] = 8'd18;
        rom[138][61] = 8'd26;
        rom[138][62] = -8'd13;
        rom[138][63] = -8'd22;
        rom[139][0] = 8'd37;
        rom[139][1] = -8'd74;
        rom[139][2] = 8'd9;
        rom[139][3] = -8'd17;
        rom[139][4] = -8'd31;
        rom[139][5] = 8'd48;
        rom[139][6] = -8'd57;
        rom[139][7] = -8'd25;
        rom[139][8] = -8'd49;
        rom[139][9] = 8'd18;
        rom[139][10] = -8'd45;
        rom[139][11] = -8'd10;
        rom[139][12] = -8'd19;
        rom[139][13] = 8'd2;
        rom[139][14] = 8'd29;
        rom[139][15] = 8'd32;
        rom[139][16] = -8'd3;
        rom[139][17] = 8'd19;
        rom[139][18] = -8'd29;
        rom[139][19] = 8'd19;
        rom[139][20] = -8'd1;
        rom[139][21] = -8'd4;
        rom[139][22] = 8'd42;
        rom[139][23] = -8'd22;
        rom[139][24] = -8'd4;
        rom[139][25] = -8'd14;
        rom[139][26] = 8'd4;
        rom[139][27] = -8'd70;
        rom[139][28] = 8'd86;
        rom[139][29] = 8'd47;
        rom[139][30] = 8'd3;
        rom[139][31] = -8'd17;
        rom[139][32] = -8'd50;
        rom[139][33] = -8'd47;
        rom[139][34] = 8'd57;
        rom[139][35] = -8'd55;
        rom[139][36] = -8'd2;
        rom[139][37] = -8'd38;
        rom[139][38] = 8'd0;
        rom[139][39] = 8'd43;
        rom[139][40] = -8'd38;
        rom[139][41] = -8'd79;
        rom[139][42] = 8'd0;
        rom[139][43] = -8'd6;
        rom[139][44] = 8'd21;
        rom[139][45] = -8'd48;
        rom[139][46] = 8'd20;
        rom[139][47] = -8'd29;
        rom[139][48] = 8'd42;
        rom[139][49] = -8'd15;
        rom[139][50] = -8'd20;
        rom[139][51] = 8'd9;
        rom[139][52] = 8'd26;
        rom[139][53] = -8'd26;
        rom[139][54] = -8'd5;
        rom[139][55] = -8'd4;
        rom[139][56] = -8'd38;
        rom[139][57] = 8'd13;
        rom[139][58] = 8'd54;
        rom[139][59] = -8'd12;
        rom[139][60] = -8'd31;
        rom[139][61] = -8'd52;
        rom[139][62] = 8'd19;
        rom[139][63] = 8'd13;
        rom[140][0] = 8'd16;
        rom[140][1] = -8'd21;
        rom[140][2] = 8'd7;
        rom[140][3] = 8'd25;
        rom[140][4] = 8'd26;
        rom[140][5] = 8'd29;
        rom[140][6] = -8'd65;
        rom[140][7] = 8'd0;
        rom[140][8] = 8'd5;
        rom[140][9] = 8'd31;
        rom[140][10] = -8'd36;
        rom[140][11] = 8'd0;
        rom[140][12] = -8'd70;
        rom[140][13] = 8'd1;
        rom[140][14] = -8'd11;
        rom[140][15] = -8'd25;
        rom[140][16] = -8'd37;
        rom[140][17] = -8'd2;
        rom[140][18] = -8'd16;
        rom[140][19] = -8'd89;
        rom[140][20] = 8'd1;
        rom[140][21] = -8'd8;
        rom[140][22] = 8'd32;
        rom[140][23] = -8'd25;
        rom[140][24] = -8'd28;
        rom[140][25] = 8'd44;
        rom[140][26] = -8'd17;
        rom[140][27] = -8'd2;
        rom[140][28] = 8'd15;
        rom[140][29] = -8'd12;
        rom[140][30] = -8'd18;
        rom[140][31] = 8'd51;
        rom[140][32] = -8'd21;
        rom[140][33] = -8'd83;
        rom[140][34] = 8'd0;
        rom[140][35] = 8'd29;
        rom[140][36] = 8'd31;
        rom[140][37] = -8'd1;
        rom[140][38] = 8'd1;
        rom[140][39] = -8'd17;
        rom[140][40] = 8'd33;
        rom[140][41] = -8'd2;
        rom[140][42] = 8'd5;
        rom[140][43] = -8'd2;
        rom[140][44] = 8'd20;
        rom[140][45] = -8'd56;
        rom[140][46] = -8'd98;
        rom[140][47] = 8'd8;
        rom[140][48] = 8'd47;
        rom[140][49] = 8'd17;
        rom[140][50] = 8'd34;
        rom[140][51] = 8'd12;
        rom[140][52] = -8'd29;
        rom[140][53] = 8'd1;
        rom[140][54] = -8'd80;
        rom[140][55] = 8'd5;
        rom[140][56] = 8'd41;
        rom[140][57] = 8'd27;
        rom[140][58] = -8'd14;
        rom[140][59] = -8'd21;
        rom[140][60] = -8'd26;
        rom[140][61] = 8'd5;
        rom[140][62] = 8'd18;
        rom[140][63] = 8'd34;
        rom[141][0] = -8'd7;
        rom[141][1] = -8'd58;
        rom[141][2] = -8'd17;
        rom[141][3] = -8'd33;
        rom[141][4] = 8'd22;
        rom[141][5] = -8'd26;
        rom[141][6] = 8'd21;
        rom[141][7] = 8'd5;
        rom[141][8] = -8'd6;
        rom[141][9] = -8'd40;
        rom[141][10] = -8'd20;
        rom[141][11] = -8'd17;
        rom[141][12] = -8'd29;
        rom[141][13] = 8'd9;
        rom[141][14] = 8'd11;
        rom[141][15] = 8'd6;
        rom[141][16] = 8'd7;
        rom[141][17] = -8'd43;
        rom[141][18] = 8'd18;
        rom[141][19] = -8'd31;
        rom[141][20] = -8'd3;
        rom[141][21] = 8'd31;
        rom[141][22] = -8'd2;
        rom[141][23] = 8'd3;
        rom[141][24] = -8'd22;
        rom[141][25] = -8'd4;
        rom[141][26] = -8'd35;
        rom[141][27] = -8'd17;
        rom[141][28] = -8'd43;
        rom[141][29] = -8'd19;
        rom[141][30] = -8'd56;
        rom[141][31] = -8'd11;
        rom[141][32] = -8'd25;
        rom[141][33] = -8'd27;
        rom[141][34] = -8'd6;
        rom[141][35] = 8'd27;
        rom[141][36] = -8'd22;
        rom[141][37] = 8'd9;
        rom[141][38] = -8'd12;
        rom[141][39] = -8'd2;
        rom[141][40] = 8'd7;
        rom[141][41] = 8'd4;
        rom[141][42] = -8'd56;
        rom[141][43] = 8'd4;
        rom[141][44] = 8'd11;
        rom[141][45] = 8'd24;
        rom[141][46] = 8'd6;
        rom[141][47] = -8'd33;
        rom[141][48] = -8'd39;
        rom[141][49] = -8'd10;
        rom[141][50] = -8'd34;
        rom[141][51] = -8'd18;
        rom[141][52] = 8'd16;
        rom[141][53] = 8'd21;
        rom[141][54] = -8'd41;
        rom[141][55] = -8'd2;
        rom[141][56] = 8'd22;
        rom[141][57] = 8'd34;
        rom[141][58] = -8'd6;
        rom[141][59] = -8'd4;
        rom[141][60] = -8'd54;
        rom[141][61] = 8'd1;
        rom[141][62] = 8'd3;
        rom[141][63] = 8'd8;
        rom[142][0] = -8'd21;
        rom[142][1] = 8'd32;
        rom[142][2] = -8'd30;
        rom[142][3] = 8'd36;
        rom[142][4] = 8'd37;
        rom[142][5] = -8'd41;
        rom[142][6] = -8'd5;
        rom[142][7] = -8'd14;
        rom[142][8] = 8'd1;
        rom[142][9] = 8'd6;
        rom[142][10] = -8'd100;
        rom[142][11] = -8'd22;
        rom[142][12] = -8'd21;
        rom[142][13] = -8'd6;
        rom[142][14] = 8'd14;
        rom[142][15] = 8'd24;
        rom[142][16] = 8'd19;
        rom[142][17] = 8'd50;
        rom[142][18] = -8'd40;
        rom[142][19] = 8'd16;
        rom[142][20] = -8'd3;
        rom[142][21] = -8'd19;
        rom[142][22] = -8'd50;
        rom[142][23] = 8'd2;
        rom[142][24] = -8'd83;
        rom[142][25] = 8'd20;
        rom[142][26] = 8'd2;
        rom[142][27] = -8'd59;
        rom[142][28] = 8'd1;
        rom[142][29] = -8'd52;
        rom[142][30] = -8'd3;
        rom[142][31] = -8'd11;
        rom[142][32] = 8'd29;
        rom[142][33] = -8'd9;
        rom[142][34] = -8'd38;
        rom[142][35] = -8'd10;
        rom[142][36] = -8'd37;
        rom[142][37] = -8'd1;
        rom[142][38] = -8'd25;
        rom[142][39] = 8'd18;
        rom[142][40] = -8'd10;
        rom[142][41] = -8'd21;
        rom[142][42] = 8'd13;
        rom[142][43] = -8'd15;
        rom[142][44] = 8'd39;
        rom[142][45] = 8'd30;
        rom[142][46] = 8'd26;
        rom[142][47] = -8'd11;
        rom[142][48] = -8'd46;
        rom[142][49] = -8'd7;
        rom[142][50] = 8'd29;
        rom[142][51] = 8'd10;
        rom[142][52] = 8'd0;
        rom[142][53] = -8'd3;
        rom[142][54] = -8'd8;
        rom[142][55] = -8'd94;
        rom[142][56] = 8'd23;
        rom[142][57] = 8'd11;
        rom[142][58] = -8'd8;
        rom[142][59] = -8'd18;
        rom[142][60] = -8'd52;
        rom[142][61] = -8'd63;
        rom[142][62] = -8'd26;
        rom[142][63] = -8'd25;
        rom[143][0] = -8'd3;
        rom[143][1] = -8'd26;
        rom[143][2] = -8'd10;
        rom[143][3] = -8'd4;
        rom[143][4] = -8'd21;
        rom[143][5] = -8'd8;
        rom[143][6] = 8'd44;
        rom[143][7] = 8'd8;
        rom[143][8] = 8'd2;
        rom[143][9] = -8'd3;
        rom[143][10] = -8'd45;
        rom[143][11] = 8'd1;
        rom[143][12] = -8'd24;
        rom[143][13] = 8'd31;
        rom[143][14] = 8'd11;
        rom[143][15] = 8'd17;
        rom[143][16] = 8'd16;
        rom[143][17] = -8'd1;
        rom[143][18] = -8'd4;
        rom[143][19] = 8'd11;
        rom[143][20] = 8'd1;
        rom[143][21] = 8'd12;
        rom[143][22] = -8'd40;
        rom[143][23] = 8'd41;
        rom[143][24] = -8'd41;
        rom[143][25] = 8'd7;
        rom[143][26] = -8'd6;
        rom[143][27] = 8'd11;
        rom[143][28] = -8'd67;
        rom[143][29] = -8'd1;
        rom[143][30] = 8'd31;
        rom[143][31] = -8'd49;
        rom[143][32] = 8'd10;
        rom[143][33] = 8'd10;
        rom[143][34] = -8'd1;
        rom[143][35] = 8'd28;
        rom[143][36] = -8'd6;
        rom[143][37] = -8'd15;
        rom[143][38] = 8'd14;
        rom[143][39] = -8'd8;
        rom[143][40] = -8'd12;
        rom[143][41] = 8'd11;
        rom[143][42] = -8'd32;
        rom[143][43] = -8'd76;
        rom[143][44] = -8'd8;
        rom[143][45] = -8'd41;
        rom[143][46] = 8'd12;
        rom[143][47] = 8'd8;
        rom[143][48] = -8'd22;
        rom[143][49] = 8'd3;
        rom[143][50] = -8'd59;
        rom[143][51] = 8'd3;
        rom[143][52] = 8'd6;
        rom[143][53] = -8'd18;
        rom[143][54] = -8'd2;
        rom[143][55] = 8'd24;
        rom[143][56] = 8'd17;
        rom[143][57] = -8'd37;
        rom[143][58] = -8'd27;
        rom[143][59] = -8'd20;
        rom[143][60] = -8'd1;
        rom[143][61] = -8'd50;
        rom[143][62] = -8'd25;
        rom[143][63] = -8'd47;
        rom[144][0] = 8'd2;
        rom[144][1] = 8'd1;
        rom[144][2] = -8'd7;
        rom[144][3] = -8'd4;
        rom[144][4] = 8'd6;
        rom[144][5] = 8'd8;
        rom[144][6] = 8'd3;
        rom[144][7] = -8'd6;
        rom[144][8] = -8'd6;
        rom[144][9] = -8'd7;
        rom[144][10] = 8'd1;
        rom[144][11] = 8'd2;
        rom[144][12] = 8'd0;
        rom[144][13] = -8'd4;
        rom[144][14] = 8'd4;
        rom[144][15] = -8'd3;
        rom[144][16] = -8'd6;
        rom[144][17] = 8'd1;
        rom[144][18] = 8'd3;
        rom[144][19] = -8'd8;
        rom[144][20] = -8'd2;
        rom[144][21] = -8'd6;
        rom[144][22] = -8'd8;
        rom[144][23] = -8'd9;
        rom[144][24] = -8'd5;
        rom[144][25] = 8'd4;
        rom[144][26] = -8'd6;
        rom[144][27] = 8'd2;
        rom[144][28] = 8'd0;
        rom[144][29] = -8'd3;
        rom[144][30] = 8'd4;
        rom[144][31] = 8'd7;
        rom[144][32] = 8'd5;
        rom[144][33] = 8'd0;
        rom[144][34] = 8'd8;
        rom[144][35] = 8'd3;
        rom[144][36] = -8'd5;
        rom[144][37] = 8'd5;
        rom[144][38] = -8'd9;
        rom[144][39] = 8'd4;
        rom[144][40] = -8'd2;
        rom[144][41] = -8'd2;
        rom[144][42] = -8'd1;
        rom[144][43] = -8'd1;
        rom[144][44] = -8'd4;
        rom[144][45] = 8'd0;
        rom[144][46] = -8'd1;
        rom[144][47] = 8'd4;
        rom[144][48] = -8'd1;
        rom[144][49] = 8'd2;
        rom[144][50] = 8'd2;
        rom[144][51] = 8'd2;
        rom[144][52] = -8'd3;
        rom[144][53] = 8'd3;
        rom[144][54] = 8'd3;
        rom[144][55] = 8'd7;
        rom[144][56] = -8'd2;
        rom[144][57] = -8'd3;
        rom[144][58] = -8'd7;
        rom[144][59] = -8'd6;
        rom[144][60] = 8'd9;
        rom[144][61] = 8'd4;
        rom[144][62] = -8'd6;
        rom[144][63] = 8'd10;
        rom[145][0] = 8'd18;
        rom[145][1] = -8'd26;
        rom[145][2] = -8'd8;
        rom[145][3] = -8'd57;
        rom[145][4] = 8'd1;
        rom[145][5] = -8'd11;
        rom[145][6] = 8'd27;
        rom[145][7] = 8'd31;
        rom[145][8] = 8'd11;
        rom[145][9] = -8'd19;
        rom[145][10] = 8'd32;
        rom[145][11] = 8'd3;
        rom[145][12] = 8'd34;
        rom[145][13] = -8'd45;
        rom[145][14] = -8'd10;
        rom[145][15] = 8'd21;
        rom[145][16] = 8'd9;
        rom[145][17] = -8'd15;
        rom[145][18] = -8'd3;
        rom[145][19] = 8'd47;
        rom[145][20] = 8'd2;
        rom[145][21] = 8'd23;
        rom[145][22] = -8'd41;
        rom[145][23] = -8'd55;
        rom[145][24] = -8'd53;
        rom[145][25] = 8'd6;
        rom[145][26] = 8'd26;
        rom[145][27] = -8'd9;
        rom[145][28] = 8'd24;
        rom[145][29] = 8'd30;
        rom[145][30] = 8'd20;
        rom[145][31] = 8'd29;
        rom[145][32] = 8'd16;
        rom[145][33] = 8'd8;
        rom[145][34] = 8'd0;
        rom[145][35] = -8'd10;
        rom[145][36] = 8'd38;
        rom[145][37] = 8'd32;
        rom[145][38] = -8'd21;
        rom[145][39] = -8'd8;
        rom[145][40] = 8'd45;
        rom[145][41] = -8'd3;
        rom[145][42] = 8'd6;
        rom[145][43] = 8'd25;
        rom[145][44] = -8'd18;
        rom[145][45] = -8'd30;
        rom[145][46] = -8'd40;
        rom[145][47] = 8'd30;
        rom[145][48] = 8'd13;
        rom[145][49] = 8'd1;
        rom[145][50] = -8'd43;
        rom[145][51] = 8'd19;
        rom[145][52] = -8'd9;
        rom[145][53] = 8'd40;
        rom[145][54] = 8'd13;
        rom[145][55] = 8'd9;
        rom[145][56] = 8'd2;
        rom[145][57] = 8'd0;
        rom[145][58] = -8'd31;
        rom[145][59] = 8'd22;
        rom[145][60] = -8'd8;
        rom[145][61] = 8'd46;
        rom[145][62] = -8'd97;
        rom[145][63] = -8'd21;
        rom[146][0] = -8'd3;
        rom[146][1] = 8'd46;
        rom[146][2] = 8'd17;
        rom[146][3] = 8'd49;
        rom[146][4] = -8'd46;
        rom[146][5] = -8'd6;
        rom[146][6] = -8'd6;
        rom[146][7] = 8'd12;
        rom[146][8] = 8'd2;
        rom[146][9] = 8'd3;
        rom[146][10] = -8'd23;
        rom[146][11] = -8'd3;
        rom[146][12] = 8'd4;
        rom[146][13] = 8'd3;
        rom[146][14] = 8'd12;
        rom[146][15] = -8'd6;
        rom[146][16] = 8'd11;
        rom[146][17] = -8'd32;
        rom[146][18] = 8'd24;
        rom[146][19] = 8'd16;
        rom[146][20] = -8'd5;
        rom[146][21] = 8'd21;
        rom[146][22] = -8'd44;
        rom[146][23] = 8'd6;
        rom[146][24] = 8'd15;
        rom[146][25] = 8'd20;
        rom[146][26] = 8'd24;
        rom[146][27] = -8'd16;
        rom[146][28] = 8'd21;
        rom[146][29] = -8'd8;
        rom[146][30] = -8'd16;
        rom[146][31] = -8'd10;
        rom[146][32] = -8'd38;
        rom[146][33] = 8'd4;
        rom[146][34] = -8'd26;
        rom[146][35] = 8'd32;
        rom[146][36] = -8'd44;
        rom[146][37] = -8'd5;
        rom[146][38] = 8'd59;
        rom[146][39] = -8'd8;
        rom[146][40] = 8'd12;
        rom[146][41] = -8'd1;
        rom[146][42] = 8'd9;
        rom[146][43] = -8'd20;
        rom[146][44] = -8'd46;
        rom[146][45] = 8'd7;
        rom[146][46] = -8'd31;
        rom[146][47] = 8'd6;
        rom[146][48] = 8'd32;
        rom[146][49] = -8'd19;
        rom[146][50] = 8'd1;
        rom[146][51] = 8'd25;
        rom[146][52] = -8'd34;
        rom[146][53] = 8'd4;
        rom[146][54] = 8'd1;
        rom[146][55] = -8'd29;
        rom[146][56] = 8'd19;
        rom[146][57] = -8'd25;
        rom[146][58] = -8'd20;
        rom[146][59] = 8'd61;
        rom[146][60] = -8'd58;
        rom[146][61] = -8'd5;
        rom[146][62] = -8'd45;
        rom[146][63] = -8'd20;
        rom[147][0] = -8'd51;
        rom[147][1] = -8'd1;
        rom[147][2] = -8'd50;
        rom[147][3] = -8'd98;
        rom[147][4] = -8'd50;
        rom[147][5] = 8'd6;
        rom[147][6] = -8'd24;
        rom[147][7] = 8'd12;
        rom[147][8] = -8'd74;
        rom[147][9] = -8'd16;
        rom[147][10] = -8'd21;
        rom[147][11] = 8'd5;
        rom[147][12] = 8'd22;
        rom[147][13] = -8'd27;
        rom[147][14] = 8'd11;
        rom[147][15] = 8'd5;
        rom[147][16] = 8'd0;
        rom[147][17] = -8'd22;
        rom[147][18] = 8'd4;
        rom[147][19] = -8'd10;
        rom[147][20] = 8'd3;
        rom[147][21] = 8'd29;
        rom[147][22] = -8'd66;
        rom[147][23] = -8'd37;
        rom[147][24] = 8'd40;
        rom[147][25] = 8'd3;
        rom[147][26] = 8'd39;
        rom[147][27] = -8'd88;
        rom[147][28] = 8'd55;
        rom[147][29] = -8'd28;
        rom[147][30] = 8'd66;
        rom[147][31] = 8'd27;
        rom[147][32] = 8'd4;
        rom[147][33] = -8'd21;
        rom[147][34] = 8'd31;
        rom[147][35] = 8'd20;
        rom[147][36] = -8'd39;
        rom[147][37] = -8'd16;
        rom[147][38] = 8'd8;
        rom[147][39] = -8'd48;
        rom[147][40] = 8'd18;
        rom[147][41] = 8'd17;
        rom[147][42] = -8'd91;
        rom[147][43] = 8'd20;
        rom[147][44] = -8'd11;
        rom[147][45] = -8'd17;
        rom[147][46] = 8'd14;
        rom[147][47] = 8'd31;
        rom[147][48] = -8'd28;
        rom[147][49] = -8'd42;
        rom[147][50] = -8'd13;
        rom[147][51] = -8'd18;
        rom[147][52] = 8'd14;
        rom[147][53] = 8'd15;
        rom[147][54] = 8'd26;
        rom[147][55] = 8'd14;
        rom[147][56] = 8'd25;
        rom[147][57] = 8'd0;
        rom[147][58] = 8'd41;
        rom[147][59] = -8'd48;
        rom[147][60] = 8'd16;
        rom[147][61] = 8'd2;
        rom[147][62] = -8'd28;
        rom[147][63] = -8'd14;
        rom[148][0] = 8'd11;
        rom[148][1] = 8'd15;
        rom[148][2] = 8'd25;
        rom[148][3] = 8'd38;
        rom[148][4] = 8'd32;
        rom[148][5] = 8'd5;
        rom[148][6] = -8'd25;
        rom[148][7] = -8'd26;
        rom[148][8] = 8'd11;
        rom[148][9] = 8'd14;
        rom[148][10] = -8'd37;
        rom[148][11] = 8'd18;
        rom[148][12] = -8'd57;
        rom[148][13] = -8'd37;
        rom[148][14] = -8'd20;
        rom[148][15] = -8'd16;
        rom[148][16] = 8'd0;
        rom[148][17] = -8'd1;
        rom[148][18] = -8'd21;
        rom[148][19] = -8'd20;
        rom[148][20] = -8'd12;
        rom[148][21] = -8'd23;
        rom[148][22] = 8'd20;
        rom[148][23] = 8'd24;
        rom[148][24] = 8'd9;
        rom[148][25] = 8'd2;
        rom[148][26] = 8'd7;
        rom[148][27] = -8'd3;
        rom[148][28] = -8'd22;
        rom[148][29] = 8'd23;
        rom[148][30] = 8'd14;
        rom[148][31] = 8'd17;
        rom[148][32] = -8'd36;
        rom[148][33] = -8'd41;
        rom[148][34] = -8'd16;
        rom[148][35] = 8'd33;
        rom[148][36] = -8'd26;
        rom[148][37] = 8'd9;
        rom[148][38] = -8'd33;
        rom[148][39] = -8'd49;
        rom[148][40] = 8'd14;
        rom[148][41] = -8'd18;
        rom[148][42] = -8'd2;
        rom[148][43] = 8'd2;
        rom[148][44] = -8'd27;
        rom[148][45] = 8'd5;
        rom[148][46] = -8'd10;
        rom[148][47] = 8'd46;
        rom[148][48] = -8'd2;
        rom[148][49] = 8'd16;
        rom[148][50] = 8'd26;
        rom[148][51] = 8'd14;
        rom[148][52] = -8'd25;
        rom[148][53] = 8'd12;
        rom[148][54] = 8'd9;
        rom[148][55] = 8'd13;
        rom[148][56] = -8'd2;
        rom[148][57] = -8'd7;
        rom[148][58] = 8'd26;
        rom[148][59] = -8'd44;
        rom[148][60] = -8'd19;
        rom[148][61] = -8'd14;
        rom[148][62] = 8'd7;
        rom[148][63] = 8'd3;
        rom[149][0] = 8'd2;
        rom[149][1] = -8'd8;
        rom[149][2] = 8'd1;
        rom[149][3] = 8'd1;
        rom[149][4] = -8'd9;
        rom[149][5] = -8'd1;
        rom[149][6] = 8'd9;
        rom[149][7] = 8'd9;
        rom[149][8] = -8'd2;
        rom[149][9] = -8'd7;
        rom[149][10] = -8'd8;
        rom[149][11] = -8'd7;
        rom[149][12] = -8'd1;
        rom[149][13] = -8'd6;
        rom[149][14] = -8'd5;
        rom[149][15] = 8'd1;
        rom[149][16] = -8'd3;
        rom[149][17] = 8'd4;
        rom[149][18] = 8'd8;
        rom[149][19] = 8'd3;
        rom[149][20] = -8'd4;
        rom[149][21] = -8'd2;
        rom[149][22] = -8'd3;
        rom[149][23] = -8'd2;
        rom[149][24] = -8'd1;
        rom[149][25] = -8'd5;
        rom[149][26] = -8'd3;
        rom[149][27] = -8'd7;
        rom[149][28] = -8'd3;
        rom[149][29] = 8'd6;
        rom[149][30] = 8'd5;
        rom[149][31] = 8'd5;
        rom[149][32] = 8'd1;
        rom[149][33] = 8'd4;
        rom[149][34] = 8'd7;
        rom[149][35] = 8'd1;
        rom[149][36] = -8'd1;
        rom[149][37] = -8'd7;
        rom[149][38] = -8'd6;
        rom[149][39] = 8'd4;
        rom[149][40] = 8'd0;
        rom[149][41] = 8'd4;
        rom[149][42] = -8'd9;
        rom[149][43] = 8'd2;
        rom[149][44] = 8'd5;
        rom[149][45] = -8'd8;
        rom[149][46] = -8'd2;
        rom[149][47] = -8'd8;
        rom[149][48] = 8'd1;
        rom[149][49] = -8'd5;
        rom[149][50] = -8'd1;
        rom[149][51] = -8'd6;
        rom[149][52] = -8'd9;
        rom[149][53] = 8'd2;
        rom[149][54] = 8'd8;
        rom[149][55] = -8'd6;
        rom[149][56] = 8'd1;
        rom[149][57] = -8'd6;
        rom[149][58] = -8'd9;
        rom[149][59] = 8'd9;
        rom[149][60] = -8'd5;
        rom[149][61] = 8'd2;
        rom[149][62] = 8'd5;
        rom[149][63] = 8'd6;
        rom[150][0] = -8'd11;
        rom[150][1] = -8'd45;
        rom[150][2] = -8'd23;
        rom[150][3] = -8'd2;
        rom[150][4] = -8'd25;
        rom[150][5] = -8'd42;
        rom[150][6] = -8'd28;
        rom[150][7] = 8'd8;
        rom[150][8] = -8'd5;
        rom[150][9] = -8'd2;
        rom[150][10] = -8'd32;
        rom[150][11] = -8'd12;
        rom[150][12] = -8'd37;
        rom[150][13] = -8'd9;
        rom[150][14] = -8'd26;
        rom[150][15] = 8'd8;
        rom[150][16] = 8'd1;
        rom[150][17] = -8'd40;
        rom[150][18] = -8'd31;
        rom[150][19] = 8'd10;
        rom[150][20] = 8'd1;
        rom[150][21] = -8'd23;
        rom[150][22] = -8'd16;
        rom[150][23] = -8'd61;
        rom[150][24] = -8'd30;
        rom[150][25] = 8'd1;
        rom[150][26] = -8'd29;
        rom[150][27] = -8'd81;
        rom[150][28] = -8'd6;
        rom[150][29] = 8'd5;
        rom[150][30] = 8'd4;
        rom[150][31] = -8'd27;
        rom[150][32] = -8'd11;
        rom[150][33] = -8'd44;
        rom[150][34] = 8'd9;
        rom[150][35] = -8'd63;
        rom[150][36] = -8'd18;
        rom[150][37] = -8'd5;
        rom[150][38] = -8'd60;
        rom[150][39] = 8'd7;
        rom[150][40] = -8'd80;
        rom[150][41] = -8'd2;
        rom[150][42] = -8'd13;
        rom[150][43] = -8'd3;
        rom[150][44] = -8'd20;
        rom[150][45] = -8'd4;
        rom[150][46] = 8'd23;
        rom[150][47] = 8'd3;
        rom[150][48] = -8'd40;
        rom[150][49] = -8'd42;
        rom[150][50] = 8'd17;
        rom[150][51] = -8'd34;
        rom[150][52] = -8'd24;
        rom[150][53] = -8'd1;
        rom[150][54] = 8'd26;
        rom[150][55] = 8'd1;
        rom[150][56] = 8'd3;
        rom[150][57] = -8'd19;
        rom[150][58] = -8'd18;
        rom[150][59] = 8'd0;
        rom[150][60] = 8'd2;
        rom[150][61] = -8'd35;
        rom[150][62] = -8'd1;
        rom[150][63] = -8'd14;
        rom[151][0] = 8'd24;
        rom[151][1] = 8'd16;
        rom[151][2] = -8'd18;
        rom[151][3] = 8'd6;
        rom[151][4] = 8'd1;
        rom[151][5] = 8'd24;
        rom[151][6] = -8'd20;
        rom[151][7] = -8'd20;
        rom[151][8] = -8'd58;
        rom[151][9] = 8'd11;
        rom[151][10] = -8'd41;
        rom[151][11] = 8'd2;
        rom[151][12] = 8'd6;
        rom[151][13] = 8'd2;
        rom[151][14] = 8'd22;
        rom[151][15] = -8'd41;
        rom[151][16] = -8'd22;
        rom[151][17] = -8'd7;
        rom[151][18] = 8'd32;
        rom[151][19] = -8'd36;
        rom[151][20] = -8'd4;
        rom[151][21] = -8'd34;
        rom[151][22] = 8'd31;
        rom[151][23] = -8'd19;
        rom[151][24] = 8'd6;
        rom[151][25] = -8'd17;
        rom[151][26] = -8'd49;
        rom[151][27] = 8'd29;
        rom[151][28] = -8'd26;
        rom[151][29] = -8'd18;
        rom[151][30] = -8'd14;
        rom[151][31] = 8'd43;
        rom[151][32] = -8'd12;
        rom[151][33] = -8'd4;
        rom[151][34] = -8'd5;
        rom[151][35] = 8'd23;
        rom[151][36] = -8'd21;
        rom[151][37] = 8'd16;
        rom[151][38] = 8'd25;
        rom[151][39] = 8'd9;
        rom[151][40] = 8'd31;
        rom[151][41] = -8'd10;
        rom[151][42] = 8'd32;
        rom[151][43] = 8'd5;
        rom[151][44] = 8'd0;
        rom[151][45] = -8'd19;
        rom[151][46] = -8'd11;
        rom[151][47] = 8'd32;
        rom[151][48] = 8'd1;
        rom[151][49] = 8'd11;
        rom[151][50] = -8'd16;
        rom[151][51] = -8'd25;
        rom[151][52] = 8'd12;
        rom[151][53] = -8'd21;
        rom[151][54] = -8'd22;
        rom[151][55] = 8'd15;
        rom[151][56] = -8'd18;
        rom[151][57] = -8'd1;
        rom[151][58] = -8'd1;
        rom[151][59] = -8'd8;
        rom[151][60] = 8'd18;
        rom[151][61] = -8'd35;
        rom[151][62] = 8'd42;
        rom[151][63] = 8'd46;
        rom[152][0] = -8'd2;
        rom[152][1] = 8'd13;
        rom[152][2] = 8'd8;
        rom[152][3] = -8'd109;
        rom[152][4] = 8'd21;
        rom[152][5] = 8'd24;
        rom[152][6] = -8'd56;
        rom[152][7] = -8'd17;
        rom[152][8] = 8'd1;
        rom[152][9] = -8'd18;
        rom[152][10] = 8'd7;
        rom[152][11] = 8'd11;
        rom[152][12] = 8'd7;
        rom[152][13] = 8'd13;
        rom[152][14] = 8'd4;
        rom[152][15] = -8'd3;
        rom[152][16] = 8'd25;
        rom[152][17] = 8'd30;
        rom[152][18] = 8'd31;
        rom[152][19] = 8'd30;
        rom[152][20] = -8'd9;
        rom[152][21] = 8'd19;
        rom[152][22] = -8'd10;
        rom[152][23] = -8'd38;
        rom[152][24] = 8'd34;
        rom[152][25] = 8'd14;
        rom[152][26] = -8'd29;
        rom[152][27] = 8'd0;
        rom[152][28] = -8'd38;
        rom[152][29] = 8'd13;
        rom[152][30] = -8'd8;
        rom[152][31] = 8'd0;
        rom[152][32] = 8'd15;
        rom[152][33] = -8'd40;
        rom[152][34] = 8'd52;
        rom[152][35] = -8'd17;
        rom[152][36] = 8'd21;
        rom[152][37] = -8'd8;
        rom[152][38] = 8'd22;
        rom[152][39] = -8'd9;
        rom[152][40] = 8'd44;
        rom[152][41] = 8'd42;
        rom[152][42] = 8'd26;
        rom[152][43] = 8'd36;
        rom[152][44] = -8'd37;
        rom[152][45] = 8'd61;
        rom[152][46] = -8'd29;
        rom[152][47] = -8'd31;
        rom[152][48] = -8'd27;
        rom[152][49] = 8'd14;
        rom[152][50] = -8'd6;
        rom[152][51] = 8'd20;
        rom[152][52] = 8'd23;
        rom[152][53] = -8'd3;
        rom[152][54] = 8'd2;
        rom[152][55] = 8'd14;
        rom[152][56] = -8'd2;
        rom[152][57] = 8'd30;
        rom[152][58] = 8'd33;
        rom[152][59] = -8'd3;
        rom[152][60] = 8'd26;
        rom[152][61] = 8'd13;
        rom[152][62] = 8'd19;
        rom[152][63] = 8'd0;
        rom[153][0] = -8'd21;
        rom[153][1] = 8'd28;
        rom[153][2] = -8'd5;
        rom[153][3] = -8'd3;
        rom[153][4] = 8'd18;
        rom[153][5] = 8'd19;
        rom[153][6] = -8'd2;
        rom[153][7] = 8'd30;
        rom[153][8] = -8'd3;
        rom[153][9] = 8'd2;
        rom[153][10] = -8'd28;
        rom[153][11] = -8'd31;
        rom[153][12] = 8'd58;
        rom[153][13] = -8'd21;
        rom[153][14] = 8'd11;
        rom[153][15] = 8'd38;
        rom[153][16] = 8'd17;
        rom[153][17] = 8'd28;
        rom[153][18] = 8'd4;
        rom[153][19] = 8'd18;
        rom[153][20] = -8'd6;
        rom[153][21] = 8'd17;
        rom[153][22] = -8'd76;
        rom[153][23] = -8'd7;
        rom[153][24] = -8'd52;
        rom[153][25] = 8'd7;
        rom[153][26] = -8'd4;
        rom[153][27] = 8'd8;
        rom[153][28] = -8'd13;
        rom[153][29] = -8'd8;
        rom[153][30] = -8'd65;
        rom[153][31] = -8'd33;
        rom[153][32] = -8'd21;
        rom[153][33] = 8'd47;
        rom[153][34] = -8'd46;
        rom[153][35] = 8'd33;
        rom[153][36] = 8'd10;
        rom[153][37] = 8'd4;
        rom[153][38] = -8'd29;
        rom[153][39] = 8'd3;
        rom[153][40] = 8'd5;
        rom[153][41] = 8'd33;
        rom[153][42] = -8'd52;
        rom[153][43] = 8'd35;
        rom[153][44] = 8'd24;
        rom[153][45] = -8'd3;
        rom[153][46] = 8'd4;
        rom[153][47] = 8'd6;
        rom[153][48] = -8'd9;
        rom[153][49] = 8'd13;
        rom[153][50] = 8'd45;
        rom[153][51] = -8'd16;
        rom[153][52] = -8'd39;
        rom[153][53] = 8'd23;
        rom[153][54] = -8'd34;
        rom[153][55] = -8'd57;
        rom[153][56] = 8'd39;
        rom[153][57] = 8'd36;
        rom[153][58] = 8'd18;
        rom[153][59] = 8'd16;
        rom[153][60] = 8'd9;
        rom[153][61] = 8'd18;
        rom[153][62] = -8'd12;
        rom[153][63] = 8'd18;
        rom[154][0] = 8'd2;
        rom[154][1] = 8'd26;
        rom[154][2] = -8'd3;
        rom[154][3] = -8'd5;
        rom[154][4] = -8'd29;
        rom[154][5] = -8'd8;
        rom[154][6] = -8'd6;
        rom[154][7] = 8'd1;
        rom[154][8] = -8'd12;
        rom[154][9] = 8'd3;
        rom[154][10] = -8'd7;
        rom[154][11] = 8'd9;
        rom[154][12] = -8'd27;
        rom[154][13] = -8'd19;
        rom[154][14] = 8'd17;
        rom[154][15] = 8'd5;
        rom[154][16] = 8'd17;
        rom[154][17] = 8'd30;
        rom[154][18] = -8'd39;
        rom[154][19] = 8'd11;
        rom[154][20] = -8'd4;
        rom[154][21] = -8'd38;
        rom[154][22] = 8'd11;
        rom[154][23] = 8'd20;
        rom[154][24] = -8'd13;
        rom[154][25] = 8'd17;
        rom[154][26] = -8'd33;
        rom[154][27] = 8'd5;
        rom[154][28] = 8'd21;
        rom[154][29] = -8'd8;
        rom[154][30] = 8'd11;
        rom[154][31] = -8'd3;
        rom[154][32] = -8'd14;
        rom[154][33] = 8'd9;
        rom[154][34] = -8'd10;
        rom[154][35] = -8'd17;
        rom[154][36] = -8'd11;
        rom[154][37] = 8'd7;
        rom[154][38] = -8'd26;
        rom[154][39] = 8'd11;
        rom[154][40] = 8'd20;
        rom[154][41] = -8'd26;
        rom[154][42] = 8'd14;
        rom[154][43] = 8'd28;
        rom[154][44] = -8'd27;
        rom[154][45] = -8'd6;
        rom[154][46] = 8'd24;
        rom[154][47] = -8'd38;
        rom[154][48] = 8'd15;
        rom[154][49] = -8'd12;
        rom[154][50] = -8'd12;
        rom[154][51] = -8'd78;
        rom[154][52] = 8'd28;
        rom[154][53] = -8'd13;
        rom[154][54] = -8'd115;
        rom[154][55] = -8'd21;
        rom[154][56] = 8'd10;
        rom[154][57] = -8'd16;
        rom[154][58] = 8'd23;
        rom[154][59] = -8'd26;
        rom[154][60] = -8'd20;
        rom[154][61] = -8'd21;
        rom[154][62] = -8'd9;
        rom[154][63] = 8'd34;
        rom[155][0] = -8'd36;
        rom[155][1] = -8'd8;
        rom[155][2] = 8'd25;
        rom[155][3] = -8'd30;
        rom[155][4] = 8'd9;
        rom[155][5] = -8'd45;
        rom[155][6] = 8'd0;
        rom[155][7] = 8'd13;
        rom[155][8] = -8'd10;
        rom[155][9] = -8'd2;
        rom[155][10] = -8'd16;
        rom[155][11] = -8'd48;
        rom[155][12] = -8'd2;
        rom[155][13] = 8'd26;
        rom[155][14] = -8'd8;
        rom[155][15] = -8'd4;
        rom[155][16] = -8'd38;
        rom[155][17] = 8'd10;
        rom[155][18] = -8'd6;
        rom[155][19] = -8'd5;
        rom[155][20] = 8'd4;
        rom[155][21] = 8'd3;
        rom[155][22] = 8'd37;
        rom[155][23] = 8'd3;
        rom[155][24] = -8'd6;
        rom[155][25] = 8'd11;
        rom[155][26] = -8'd3;
        rom[155][27] = -8'd5;
        rom[155][28] = 8'd21;
        rom[155][29] = 8'd1;
        rom[155][30] = -8'd40;
        rom[155][31] = -8'd4;
        rom[155][32] = -8'd23;
        rom[155][33] = -8'd10;
        rom[155][34] = 8'd30;
        rom[155][35] = 8'd35;
        rom[155][36] = -8'd15;
        rom[155][37] = 8'd0;
        rom[155][38] = 8'd16;
        rom[155][39] = -8'd3;
        rom[155][40] = 8'd26;
        rom[155][41] = 8'd36;
        rom[155][42] = -8'd36;
        rom[155][43] = 8'd10;
        rom[155][44] = -8'd25;
        rom[155][45] = -8'd10;
        rom[155][46] = -8'd13;
        rom[155][47] = 8'd49;
        rom[155][48] = 8'd31;
        rom[155][49] = -8'd14;
        rom[155][50] = 8'd37;
        rom[155][51] = 8'd7;
        rom[155][52] = -8'd1;
        rom[155][53] = 8'd18;
        rom[155][54] = 8'd39;
        rom[155][55] = -8'd1;
        rom[155][56] = 8'd59;
        rom[155][57] = 8'd22;
        rom[155][58] = -8'd3;
        rom[155][59] = -8'd6;
        rom[155][60] = 8'd29;
        rom[155][61] = 8'd23;
        rom[155][62] = -8'd10;
        rom[155][63] = -8'd38;
        rom[156][0] = 8'd7;
        rom[156][1] = 8'd28;
        rom[156][2] = 8'd24;
        rom[156][3] = -8'd23;
        rom[156][4] = 8'd26;
        rom[156][5] = -8'd5;
        rom[156][6] = 8'd33;
        rom[156][7] = 8'd39;
        rom[156][8] = -8'd42;
        rom[156][9] = 8'd5;
        rom[156][10] = -8'd73;
        rom[156][11] = -8'd1;
        rom[156][12] = -8'd37;
        rom[156][13] = -8'd35;
        rom[156][14] = 8'd38;
        rom[156][15] = -8'd16;
        rom[156][16] = -8'd81;
        rom[156][17] = 8'd6;
        rom[156][18] = -8'd99;
        rom[156][19] = 8'd33;
        rom[156][20] = -8'd13;
        rom[156][21] = 8'd10;
        rom[156][22] = 8'd30;
        rom[156][23] = -8'd13;
        rom[156][24] = -8'd10;
        rom[156][25] = -8'd22;
        rom[156][26] = 8'd15;
        rom[156][27] = 8'd26;
        rom[156][28] = -8'd10;
        rom[156][29] = 8'd28;
        rom[156][30] = -8'd29;
        rom[156][31] = 8'd5;
        rom[156][32] = -8'd13;
        rom[156][33] = -8'd42;
        rom[156][34] = -8'd40;
        rom[156][35] = 8'd25;
        rom[156][36] = -8'd1;
        rom[156][37] = -8'd23;
        rom[156][38] = 8'd37;
        rom[156][39] = 8'd35;
        rom[156][40] = -8'd47;
        rom[156][41] = 8'd32;
        rom[156][42] = 8'd23;
        rom[156][43] = 8'd52;
        rom[156][44] = -8'd10;
        rom[156][45] = -8'd2;
        rom[156][46] = -8'd9;
        rom[156][47] = 8'd24;
        rom[156][48] = -8'd3;
        rom[156][49] = -8'd16;
        rom[156][50] = 8'd4;
        rom[156][51] = 8'd35;
        rom[156][52] = -8'd8;
        rom[156][53] = 8'd9;
        rom[156][54] = -8'd23;
        rom[156][55] = -8'd16;
        rom[156][56] = 8'd30;
        rom[156][57] = 8'd45;
        rom[156][58] = 8'd37;
        rom[156][59] = 8'd19;
        rom[156][60] = 8'd19;
        rom[156][61] = 8'd21;
        rom[156][62] = -8'd32;
        rom[156][63] = 8'd31;
        rom[157][0] = -8'd64;
        rom[157][1] = 8'd16;
        rom[157][2] = -8'd59;
        rom[157][3] = -8'd32;
        rom[157][4] = -8'd48;
        rom[157][5] = 8'd5;
        rom[157][6] = -8'd16;
        rom[157][7] = -8'd21;
        rom[157][8] = 8'd4;
        rom[157][9] = -8'd3;
        rom[157][10] = -8'd18;
        rom[157][11] = 8'd20;
        rom[157][12] = -8'd16;
        rom[157][13] = -8'd15;
        rom[157][14] = 8'd26;
        rom[157][15] = -8'd52;
        rom[157][16] = -8'd8;
        rom[157][17] = 8'd28;
        rom[157][18] = -8'd6;
        rom[157][19] = -8'd43;
        rom[157][20] = -8'd5;
        rom[157][21] = 8'd14;
        rom[157][22] = 8'd21;
        rom[157][23] = -8'd93;
        rom[157][24] = 8'd14;
        rom[157][25] = -8'd20;
        rom[157][26] = 8'd32;
        rom[157][27] = -8'd9;
        rom[157][28] = 8'd25;
        rom[157][29] = 8'd10;
        rom[157][30] = -8'd76;
        rom[157][31] = 8'd10;
        rom[157][32] = -8'd21;
        rom[157][33] = -8'd43;
        rom[157][34] = 8'd6;
        rom[157][35] = 8'd29;
        rom[157][36] = -8'd5;
        rom[157][37] = -8'd1;
        rom[157][38] = -8'd17;
        rom[157][39] = -8'd94;
        rom[157][40] = -8'd6;
        rom[157][41] = 8'd2;
        rom[157][42] = 8'd10;
        rom[157][43] = -8'd39;
        rom[157][44] = 8'd4;
        rom[157][45] = 8'd9;
        rom[157][46] = -8'd52;
        rom[157][47] = 8'd0;
        rom[157][48] = -8'd1;
        rom[157][49] = -8'd33;
        rom[157][50] = 8'd5;
        rom[157][51] = 8'd29;
        rom[157][52] = -8'd46;
        rom[157][53] = -8'd11;
        rom[157][54] = 8'd6;
        rom[157][55] = -8'd45;
        rom[157][56] = -8'd64;
        rom[157][57] = -8'd9;
        rom[157][58] = -8'd48;
        rom[157][59] = -8'd80;
        rom[157][60] = 8'd11;
        rom[157][61] = 8'd21;
        rom[157][62] = -8'd16;
        rom[157][63] = -8'd8;
        rom[158][0] = -8'd16;
        rom[158][1] = 8'd18;
        rom[158][2] = -8'd19;
        rom[158][3] = 8'd25;
        rom[158][4] = -8'd29;
        rom[158][5] = -8'd37;
        rom[158][6] = 8'd21;
        rom[158][7] = 8'd14;
        rom[158][8] = 8'd10;
        rom[158][9] = 8'd14;
        rom[158][10] = 8'd5;
        rom[158][11] = -8'd3;
        rom[158][12] = -8'd52;
        rom[158][13] = 8'd19;
        rom[158][14] = -8'd14;
        rom[158][15] = -8'd17;
        rom[158][16] = 8'd3;
        rom[158][17] = -8'd7;
        rom[158][18] = 8'd31;
        rom[158][19] = -8'd5;
        rom[158][20] = -8'd6;
        rom[158][21] = -8'd8;
        rom[158][22] = -8'd17;
        rom[158][23] = -8'd9;
        rom[158][24] = 8'd15;
        rom[158][25] = 8'd30;
        rom[158][26] = -8'd17;
        rom[158][27] = -8'd9;
        rom[158][28] = -8'd7;
        rom[158][29] = 8'd17;
        rom[158][30] = -8'd23;
        rom[158][31] = -8'd18;
        rom[158][32] = -8'd6;
        rom[158][33] = -8'd27;
        rom[158][34] = 8'd9;
        rom[158][35] = 8'd16;
        rom[158][36] = 8'd28;
        rom[158][37] = 8'd31;
        rom[158][38] = 8'd0;
        rom[158][39] = 8'd14;
        rom[158][40] = 8'd32;
        rom[158][41] = -8'd26;
        rom[158][42] = -8'd4;
        rom[158][43] = -8'd7;
        rom[158][44] = -8'd55;
        rom[158][45] = 8'd23;
        rom[158][46] = 8'd3;
        rom[158][47] = 8'd10;
        rom[158][48] = 8'd12;
        rom[158][49] = 8'd6;
        rom[158][50] = -8'd96;
        rom[158][51] = -8'd47;
        rom[158][52] = 8'd12;
        rom[158][53] = -8'd6;
        rom[158][54] = -8'd37;
        rom[158][55] = 8'd18;
        rom[158][56] = 8'd4;
        rom[158][57] = -8'd11;
        rom[158][58] = -8'd49;
        rom[158][59] = -8'd10;
        rom[158][60] = -8'd52;
        rom[158][61] = 8'd7;
        rom[158][62] = 8'd16;
        rom[158][63] = 8'd8;
        rom[159][0] = 8'd36;
        rom[159][1] = -8'd2;
        rom[159][2] = 8'd17;
        rom[159][3] = -8'd46;
        rom[159][4] = -8'd30;
        rom[159][5] = -8'd41;
        rom[159][6] = 8'd54;
        rom[159][7] = 8'd36;
        rom[159][8] = -8'd3;
        rom[159][9] = -8'd13;
        rom[159][10] = -8'd15;
        rom[159][11] = -8'd13;
        rom[159][12] = 8'd5;
        rom[159][13] = -8'd20;
        rom[159][14] = 8'd7;
        rom[159][15] = 8'd27;
        rom[159][16] = -8'd6;
        rom[159][17] = 8'd10;
        rom[159][18] = -8'd3;
        rom[159][19] = 8'd28;
        rom[159][20] = 8'd4;
        rom[159][21] = 8'd2;
        rom[159][22] = 8'd7;
        rom[159][23] = -8'd3;
        rom[159][24] = 8'd9;
        rom[159][25] = -8'd3;
        rom[159][26] = 8'd1;
        rom[159][27] = -8'd20;
        rom[159][28] = -8'd25;
        rom[159][29] = 8'd23;
        rom[159][30] = -8'd12;
        rom[159][31] = 8'd46;
        rom[159][32] = 8'd39;
        rom[159][33] = -8'd24;
        rom[159][34] = -8'd8;
        rom[159][35] = -8'd12;
        rom[159][36] = 8'd35;
        rom[159][37] = 8'd49;
        rom[159][38] = 8'd23;
        rom[159][39] = 8'd12;
        rom[159][40] = -8'd13;
        rom[159][41] = 8'd30;
        rom[159][42] = -8'd16;
        rom[159][43] = 8'd2;
        rom[159][44] = 8'd5;
        rom[159][45] = -8'd19;
        rom[159][46] = -8'd14;
        rom[159][47] = -8'd8;
        rom[159][48] = -8'd41;
        rom[159][49] = 8'd25;
        rom[159][50] = 8'd9;
        rom[159][51] = -8'd6;
        rom[159][52] = -8'd34;
        rom[159][53] = -8'd20;
        rom[159][54] = -8'd28;
        rom[159][55] = 8'd12;
        rom[159][56] = -8'd69;
        rom[159][57] = 8'd0;
        rom[159][58] = 8'd33;
        rom[159][59] = -8'd31;
        rom[159][60] = 8'd52;
        rom[159][61] = 8'd50;
        rom[159][62] = 8'd0;
        rom[159][63] = -8'd19;
        rom[160][0] = 8'd3;
        rom[160][1] = 8'd11;
        rom[160][2] = -8'd15;
        rom[160][3] = 8'd9;
        rom[160][4] = 8'd7;
        rom[160][5] = -8'd23;
        rom[160][6] = -8'd33;
        rom[160][7] = 8'd3;
        rom[160][8] = -8'd12;
        rom[160][9] = -8'd10;
        rom[160][10] = -8'd37;
        rom[160][11] = -8'd54;
        rom[160][12] = -8'd2;
        rom[160][13] = 8'd14;
        rom[160][14] = 8'd8;
        rom[160][15] = -8'd31;
        rom[160][16] = -8'd10;
        rom[160][17] = 8'd12;
        rom[160][18] = 8'd48;
        rom[160][19] = 8'd12;
        rom[160][20] = 8'd0;
        rom[160][21] = 8'd8;
        rom[160][22] = 8'd0;
        rom[160][23] = 8'd20;
        rom[160][24] = -8'd98;
        rom[160][25] = -8'd1;
        rom[160][26] = 8'd38;
        rom[160][27] = 8'd0;
        rom[160][28] = 8'd19;
        rom[160][29] = -8'd28;
        rom[160][30] = -8'd44;
        rom[160][31] = -8'd21;
        rom[160][32] = 8'd31;
        rom[160][33] = 8'd60;
        rom[160][34] = -8'd52;
        rom[160][35] = -8'd6;
        rom[160][36] = 8'd5;
        rom[160][37] = 8'd44;
        rom[160][38] = 8'd43;
        rom[160][39] = -8'd36;
        rom[160][40] = 8'd7;
        rom[160][41] = 8'd32;
        rom[160][42] = 8'd29;
        rom[160][43] = -8'd49;
        rom[160][44] = 8'd10;
        rom[160][45] = 8'd15;
        rom[160][46] = 8'd2;
        rom[160][47] = 8'd33;
        rom[160][48] = -8'd13;
        rom[160][49] = -8'd19;
        rom[160][50] = -8'd16;
        rom[160][51] = -8'd24;
        rom[160][52] = 8'd9;
        rom[160][53] = -8'd18;
        rom[160][54] = -8'd18;
        rom[160][55] = -8'd23;
        rom[160][56] = -8'd9;
        rom[160][57] = 8'd6;
        rom[160][58] = -8'd18;
        rom[160][59] = -8'd21;
        rom[160][60] = -8'd43;
        rom[160][61] = -8'd17;
        rom[160][62] = 8'd9;
        rom[160][63] = -8'd30;
        rom[161][0] = -8'd22;
        rom[161][1] = 8'd19;
        rom[161][2] = -8'd16;
        rom[161][3] = -8'd17;
        rom[161][4] = -8'd31;
        rom[161][5] = 8'd18;
        rom[161][6] = -8'd55;
        rom[161][7] = 8'd12;
        rom[161][8] = 8'd13;
        rom[161][9] = -8'd40;
        rom[161][10] = -8'd4;
        rom[161][11] = -8'd3;
        rom[161][12] = 8'd11;
        rom[161][13] = -8'd76;
        rom[161][14] = 8'd49;
        rom[161][15] = 8'd6;
        rom[161][16] = 8'd10;
        rom[161][17] = 8'd40;
        rom[161][18] = 8'd24;
        rom[161][19] = -8'd40;
        rom[161][20] = -8'd8;
        rom[161][21] = -8'd14;
        rom[161][22] = -8'd21;
        rom[161][23] = -8'd76;
        rom[161][24] = 8'd18;
        rom[161][25] = -8'd13;
        rom[161][26] = -8'd1;
        rom[161][27] = -8'd18;
        rom[161][28] = -8'd9;
        rom[161][29] = -8'd28;
        rom[161][30] = -8'd21;
        rom[161][31] = 8'd19;
        rom[161][32] = -8'd36;
        rom[161][33] = 8'd28;
        rom[161][34] = -8'd11;
        rom[161][35] = 8'd9;
        rom[161][36] = -8'd1;
        rom[161][37] = 8'd14;
        rom[161][38] = -8'd34;
        rom[161][39] = 8'd12;
        rom[161][40] = -8'd31;
        rom[161][41] = -8'd13;
        rom[161][42] = -8'd26;
        rom[161][43] = -8'd13;
        rom[161][44] = 8'd7;
        rom[161][45] = 8'd4;
        rom[161][46] = -8'd19;
        rom[161][47] = -8'd14;
        rom[161][48] = 8'd41;
        rom[161][49] = 8'd26;
        rom[161][50] = 8'd19;
        rom[161][51] = -8'd20;
        rom[161][52] = -8'd92;
        rom[161][53] = -8'd38;
        rom[161][54] = -8'd39;
        rom[161][55] = -8'd20;
        rom[161][56] = -8'd24;
        rom[161][57] = -8'd21;
        rom[161][58] = -8'd23;
        rom[161][59] = -8'd16;
        rom[161][60] = -8'd42;
        rom[161][61] = 8'd16;
        rom[161][62] = 8'd29;
        rom[161][63] = -8'd23;
        rom[162][0] = -8'd12;
        rom[162][1] = 8'd26;
        rom[162][2] = -8'd48;
        rom[162][3] = -8'd17;
        rom[162][4] = -8'd4;
        rom[162][5] = 8'd10;
        rom[162][6] = -8'd59;
        rom[162][7] = 8'd14;
        rom[162][8] = 8'd48;
        rom[162][9] = -8'd10;
        rom[162][10] = 8'd3;
        rom[162][11] = 8'd23;
        rom[162][12] = -8'd20;
        rom[162][13] = 8'd19;
        rom[162][14] = -8'd26;
        rom[162][15] = -8'd22;
        rom[162][16] = 8'd11;
        rom[162][17] = -8'd30;
        rom[162][18] = 8'd14;
        rom[162][19] = 8'd44;
        rom[162][20] = -8'd6;
        rom[162][21] = 8'd2;
        rom[162][22] = 8'd16;
        rom[162][23] = 8'd6;
        rom[162][24] = 8'd16;
        rom[162][25] = 8'd20;
        rom[162][26] = 8'd8;
        rom[162][27] = -8'd65;
        rom[162][28] = -8'd13;
        rom[162][29] = -8'd77;
        rom[162][30] = -8'd39;
        rom[162][31] = 8'd1;
        rom[162][32] = -8'd1;
        rom[162][33] = 8'd18;
        rom[162][34] = 8'd26;
        rom[162][35] = -8'd40;
        rom[162][36] = -8'd19;
        rom[162][37] = -8'd24;
        rom[162][38] = 8'd10;
        rom[162][39] = 8'd6;
        rom[162][40] = 8'd9;
        rom[162][41] = -8'd30;
        rom[162][42] = -8'd23;
        rom[162][43] = -8'd36;
        rom[162][44] = -8'd50;
        rom[162][45] = -8'd10;
        rom[162][46] = 8'd26;
        rom[162][47] = -8'd54;
        rom[162][48] = -8'd18;
        rom[162][49] = 8'd25;
        rom[162][50] = -8'd29;
        rom[162][51] = 8'd23;
        rom[162][52] = -8'd17;
        rom[162][53] = 8'd5;
        rom[162][54] = -8'd7;
        rom[162][55] = -8'd25;
        rom[162][56] = -8'd9;
        rom[162][57] = 8'd3;
        rom[162][58] = -8'd13;
        rom[162][59] = -8'd46;
        rom[162][60] = -8'd64;
        rom[162][61] = -8'd29;
        rom[162][62] = -8'd5;
        rom[162][63] = -8'd34;
        rom[163][0] = -8'd46;
        rom[163][1] = 8'd18;
        rom[163][2] = 8'd25;
        rom[163][3] = 8'd66;
        rom[163][4] = 8'd10;
        rom[163][5] = -8'd4;
        rom[163][6] = -8'd77;
        rom[163][7] = -8'd34;
        rom[163][8] = 8'd2;
        rom[163][9] = -8'd57;
        rom[163][10] = -8'd29;
        rom[163][11] = 8'd20;
        rom[163][12] = 8'd16;
        rom[163][13] = -8'd10;
        rom[163][14] = -8'd20;
        rom[163][15] = -8'd4;
        rom[163][16] = 8'd1;
        rom[163][17] = 8'd9;
        rom[163][18] = -8'd29;
        rom[163][19] = -8'd18;
        rom[163][20] = -8'd11;
        rom[163][21] = 8'd23;
        rom[163][22] = -8'd19;
        rom[163][23] = -8'd35;
        rom[163][24] = -8'd5;
        rom[163][25] = -8'd41;
        rom[163][26] = -8'd42;
        rom[163][27] = -8'd5;
        rom[163][28] = -8'd2;
        rom[163][29] = -8'd44;
        rom[163][30] = 8'd31;
        rom[163][31] = -8'd21;
        rom[163][32] = -8'd56;
        rom[163][33] = -8'd49;
        rom[163][34] = 8'd25;
        rom[163][35] = -8'd2;
        rom[163][36] = -8'd22;
        rom[163][37] = -8'd11;
        rom[163][38] = -8'd63;
        rom[163][39] = 8'd31;
        rom[163][40] = -8'd8;
        rom[163][41] = -8'd22;
        rom[163][42] = 8'd0;
        rom[163][43] = 8'd35;
        rom[163][44] = 8'd3;
        rom[163][45] = 8'd9;
        rom[163][46] = -8'd2;
        rom[163][47] = -8'd6;
        rom[163][48] = 8'd48;
        rom[163][49] = 8'd9;
        rom[163][50] = 8'd9;
        rom[163][51] = 8'd26;
        rom[163][52] = 8'd24;
        rom[163][53] = -8'd40;
        rom[163][54] = -8'd31;
        rom[163][55] = -8'd44;
        rom[163][56] = 8'd49;
        rom[163][57] = 8'd30;
        rom[163][58] = 8'd4;
        rom[163][59] = 8'd24;
        rom[163][60] = -8'd31;
        rom[163][61] = -8'd28;
        rom[163][62] = -8'd35;
        rom[163][63] = 8'd38;
        rom[164][0] = 8'd21;
        rom[164][1] = 8'd4;
        rom[164][2] = 8'd27;
        rom[164][3] = 8'd21;
        rom[164][4] = 8'd21;
        rom[164][5] = 8'd11;
        rom[164][6] = -8'd79;
        rom[164][7] = 8'd15;
        rom[164][8] = 8'd37;
        rom[164][9] = -8'd13;
        rom[164][10] = -8'd23;
        rom[164][11] = -8'd8;
        rom[164][12] = -8'd27;
        rom[164][13] = -8'd38;
        rom[164][14] = -8'd23;
        rom[164][15] = -8'd29;
        rom[164][16] = 8'd18;
        rom[164][17] = -8'd2;
        rom[164][18] = 8'd2;
        rom[164][19] = -8'd4;
        rom[164][20] = -8'd2;
        rom[164][21] = 8'd16;
        rom[164][22] = -8'd8;
        rom[164][23] = -8'd25;
        rom[164][24] = -8'd23;
        rom[164][25] = 8'd4;
        rom[164][26] = -8'd6;
        rom[164][27] = -8'd24;
        rom[164][28] = 8'd33;
        rom[164][29] = -8'd3;
        rom[164][30] = -8'd10;
        rom[164][31] = 8'd2;
        rom[164][32] = -8'd80;
        rom[164][33] = -8'd24;
        rom[164][34] = -8'd6;
        rom[164][35] = -8'd17;
        rom[164][36] = 8'd14;
        rom[164][37] = 8'd17;
        rom[164][38] = 8'd9;
        rom[164][39] = 8'd10;
        rom[164][40] = -8'd4;
        rom[164][41] = -8'd31;
        rom[164][42] = -8'd11;
        rom[164][43] = 8'd18;
        rom[164][44] = -8'd58;
        rom[164][45] = -8'd5;
        rom[164][46] = -8'd62;
        rom[164][47] = -8'd8;
        rom[164][48] = -8'd4;
        rom[164][49] = -8'd8;
        rom[164][50] = 8'd9;
        rom[164][51] = -8'd24;
        rom[164][52] = -8'd40;
        rom[164][53] = 8'd53;
        rom[164][54] = 8'd0;
        rom[164][55] = 8'd12;
        rom[164][56] = -8'd30;
        rom[164][57] = 8'd25;
        rom[164][58] = -8'd24;
        rom[164][59] = 8'd47;
        rom[164][60] = -8'd31;
        rom[164][61] = -8'd5;
        rom[164][62] = -8'd17;
        rom[164][63] = -8'd24;
        rom[165][0] = -8'd38;
        rom[165][1] = -8'd29;
        rom[165][2] = -8'd15;
        rom[165][3] = -8'd86;
        rom[165][4] = -8'd23;
        rom[165][5] = -8'd32;
        rom[165][6] = -8'd47;
        rom[165][7] = -8'd18;
        rom[165][8] = 8'd10;
        rom[165][9] = 8'd28;
        rom[165][10] = -8'd73;
        rom[165][11] = -8'd45;
        rom[165][12] = -8'd35;
        rom[165][13] = 8'd32;
        rom[165][14] = 8'd30;
        rom[165][15] = 8'd5;
        rom[165][16] = -8'd34;
        rom[165][17] = 8'd29;
        rom[165][18] = 8'd16;
        rom[165][19] = -8'd79;
        rom[165][20] = -8'd1;
        rom[165][21] = -8'd22;
        rom[165][22] = -8'd35;
        rom[165][23] = -8'd31;
        rom[165][24] = -8'd9;
        rom[165][25] = 8'd8;
        rom[165][26] = 8'd3;
        rom[165][27] = -8'd41;
        rom[165][28] = 8'd4;
        rom[165][29] = 8'd4;
        rom[165][30] = -8'd65;
        rom[165][31] = -8'd17;
        rom[165][32] = -8'd92;
        rom[165][33] = 8'd41;
        rom[165][34] = -8'd51;
        rom[165][35] = -8'd10;
        rom[165][36] = 8'd12;
        rom[165][37] = -8'd33;
        rom[165][38] = -8'd38;
        rom[165][39] = 8'd13;
        rom[165][40] = 8'd53;
        rom[165][41] = 8'd3;
        rom[165][42] = -8'd12;
        rom[165][43] = 8'd19;
        rom[165][44] = -8'd100;
        rom[165][45] = -8'd21;
        rom[165][46] = 8'd7;
        rom[165][47] = -8'd20;
        rom[165][48] = -8'd23;
        rom[165][49] = 8'd40;
        rom[165][50] = 8'd15;
        rom[165][51] = -8'd6;
        rom[165][52] = 8'd12;
        rom[165][53] = 8'd9;
        rom[165][54] = -8'd43;
        rom[165][55] = -8'd10;
        rom[165][56] = -8'd52;
        rom[165][57] = 8'd22;
        rom[165][58] = -8'd3;
        rom[165][59] = -8'd22;
        rom[165][60] = -8'd4;
        rom[165][61] = 8'd5;
        rom[165][62] = -8'd3;
        rom[165][63] = -8'd67;
        rom[166][0] = 8'd25;
        rom[166][1] = 8'd13;
        rom[166][2] = 8'd23;
        rom[166][3] = -8'd2;
        rom[166][4] = -8'd27;
        rom[166][5] = 8'd3;
        rom[166][6] = 8'd32;
        rom[166][7] = 8'd61;
        rom[166][8] = 8'd0;
        rom[166][9] = 8'd56;
        rom[166][10] = -8'd39;
        rom[166][11] = 8'd0;
        rom[166][12] = -8'd11;
        rom[166][13] = -8'd28;
        rom[166][14] = -8'd11;
        rom[166][15] = 8'd33;
        rom[166][16] = 8'd45;
        rom[166][17] = -8'd2;
        rom[166][18] = 8'd7;
        rom[166][19] = 8'd2;
        rom[166][20] = -8'd6;
        rom[166][21] = -8'd21;
        rom[166][22] = -8'd38;
        rom[166][23] = -8'd17;
        rom[166][24] = 8'd9;
        rom[166][25] = 8'd24;
        rom[166][26] = 8'd41;
        rom[166][27] = 8'd21;
        rom[166][28] = 8'd17;
        rom[166][29] = 8'd31;
        rom[166][30] = -8'd1;
        rom[166][31] = 8'd50;
        rom[166][32] = -8'd7;
        rom[166][33] = -8'd8;
        rom[166][34] = -8'd4;
        rom[166][35] = 8'd36;
        rom[166][36] = 8'd26;
        rom[166][37] = 8'd1;
        rom[166][38] = -8'd37;
        rom[166][39] = -8'd54;
        rom[166][40] = -8'd15;
        rom[166][41] = -8'd59;
        rom[166][42] = -8'd28;
        rom[166][43] = 8'd42;
        rom[166][44] = 8'd44;
        rom[166][45] = -8'd21;
        rom[166][46] = -8'd21;
        rom[166][47] = -8'd15;
        rom[166][48] = -8'd1;
        rom[166][49] = -8'd10;
        rom[166][50] = -8'd26;
        rom[166][51] = -8'd1;
        rom[166][52] = 8'd16;
        rom[166][53] = 8'd56;
        rom[166][54] = 8'd17;
        rom[166][55] = 8'd28;
        rom[166][56] = -8'd64;
        rom[166][57] = -8'd27;
        rom[166][58] = -8'd29;
        rom[166][59] = 8'd34;
        rom[166][60] = 8'd24;
        rom[166][61] = -8'd21;
        rom[166][62] = -8'd32;
        rom[166][63] = -8'd28;
        rom[167][0] = 8'd22;
        rom[167][1] = 8'd22;
        rom[167][2] = -8'd3;
        rom[167][3] = 8'd34;
        rom[167][4] = -8'd32;
        rom[167][5] = 8'd13;
        rom[167][6] = 8'd15;
        rom[167][7] = 8'd24;
        rom[167][8] = 8'd73;
        rom[167][9] = 8'd3;
        rom[167][10] = -8'd28;
        rom[167][11] = 8'd47;
        rom[167][12] = -8'd56;
        rom[167][13] = 8'd24;
        rom[167][14] = 8'd31;
        rom[167][15] = 8'd39;
        rom[167][16] = 8'd14;
        rom[167][17] = -8'd8;
        rom[167][18] = 8'd42;
        rom[167][19] = 8'd28;
        rom[167][20] = 8'd0;
        rom[167][21] = 8'd0;
        rom[167][22] = -8'd11;
        rom[167][23] = 8'd20;
        rom[167][24] = 8'd51;
        rom[167][25] = -8'd45;
        rom[167][26] = 8'd15;
        rom[167][27] = 8'd17;
        rom[167][28] = 8'd8;
        rom[167][29] = 8'd44;
        rom[167][30] = -8'd31;
        rom[167][31] = -8'd11;
        rom[167][32] = -8'd13;
        rom[167][33] = -8'd69;
        rom[167][34] = -8'd17;
        rom[167][35] = 8'd23;
        rom[167][36] = 8'd7;
        rom[167][37] = -8'd23;
        rom[167][38] = 8'd7;
        rom[167][39] = 8'd35;
        rom[167][40] = -8'd7;
        rom[167][41] = -8'd21;
        rom[167][42] = 8'd16;
        rom[167][43] = -8'd21;
        rom[167][44] = -8'd45;
        rom[167][45] = 8'd23;
        rom[167][46] = 8'd20;
        rom[167][47] = -8'd23;
        rom[167][48] = 8'd33;
        rom[167][49] = 8'd4;
        rom[167][50] = -8'd1;
        rom[167][51] = 8'd35;
        rom[167][52] = -8'd10;
        rom[167][53] = -8'd8;
        rom[167][54] = 8'd24;
        rom[167][55] = -8'd44;
        rom[167][56] = -8'd21;
        rom[167][57] = 8'd2;
        rom[167][58] = -8'd17;
        rom[167][59] = 8'd6;
        rom[167][60] = 8'd6;
        rom[167][61] = 8'd1;
        rom[167][62] = 8'd6;
        rom[167][63] = 8'd25;
        rom[168][0] = -8'd31;
        rom[168][1] = -8'd16;
        rom[168][2] = -8'd29;
        rom[168][3] = 8'd15;
        rom[168][4] = -8'd33;
        rom[168][5] = 8'd17;
        rom[168][6] = 8'd29;
        rom[168][7] = -8'd10;
        rom[168][8] = -8'd14;
        rom[168][9] = -8'd18;
        rom[168][10] = -8'd16;
        rom[168][11] = -8'd5;
        rom[168][12] = 8'd22;
        rom[168][13] = 8'd33;
        rom[168][14] = -8'd62;
        rom[168][15] = -8'd32;
        rom[168][16] = -8'd7;
        rom[168][17] = -8'd16;
        rom[168][18] = -8'd8;
        rom[168][19] = -8'd34;
        rom[168][20] = -8'd11;
        rom[168][21] = 8'd22;
        rom[168][22] = -8'd18;
        rom[168][23] = 8'd12;
        rom[168][24] = -8'd20;
        rom[168][25] = -8'd26;
        rom[168][26] = 8'd19;
        rom[168][27] = 8'd26;
        rom[168][28] = 8'd37;
        rom[168][29] = -8'd128;
        rom[168][30] = 8'd19;
        rom[168][31] = 8'd31;
        rom[168][32] = -8'd28;
        rom[168][33] = -8'd19;
        rom[168][34] = -8'd10;
        rom[168][35] = -8'd8;
        rom[168][36] = -8'd30;
        rom[168][37] = -8'd2;
        rom[168][38] = -8'd12;
        rom[168][39] = -8'd15;
        rom[168][40] = 8'd21;
        rom[168][41] = -8'd15;
        rom[168][42] = -8'd32;
        rom[168][43] = 8'd12;
        rom[168][44] = 8'd17;
        rom[168][45] = -8'd50;
        rom[168][46] = 8'd20;
        rom[168][47] = -8'd24;
        rom[168][48] = -8'd20;
        rom[168][49] = 8'd3;
        rom[168][50] = -8'd29;
        rom[168][51] = -8'd18;
        rom[168][52] = -8'd27;
        rom[168][53] = 8'd12;
        rom[168][54] = 8'd2;
        rom[168][55] = -8'd35;
        rom[168][56] = 8'd6;
        rom[168][57] = 8'd21;
        rom[168][58] = -8'd46;
        rom[168][59] = 8'd39;
        rom[168][60] = -8'd19;
        rom[168][61] = -8'd20;
        rom[168][62] = -8'd50;
        rom[168][63] = 8'd21;
        rom[169][0] = 8'd13;
        rom[169][1] = 8'd1;
        rom[169][2] = 8'd17;
        rom[169][3] = 8'd23;
        rom[169][4] = 8'd29;
        rom[169][5] = 8'd14;
        rom[169][6] = 8'd8;
        rom[169][7] = 8'd10;
        rom[169][8] = 8'd21;
        rom[169][9] = 8'd18;
        rom[169][10] = -8'd61;
        rom[169][11] = 8'd46;
        rom[169][12] = -8'd16;
        rom[169][13] = -8'd13;
        rom[169][14] = 8'd5;
        rom[169][15] = 8'd29;
        rom[169][16] = -8'd17;
        rom[169][17] = -8'd36;
        rom[169][18] = -8'd29;
        rom[169][19] = 8'd12;
        rom[169][20] = -8'd10;
        rom[169][21] = 8'd12;
        rom[169][22] = 8'd8;
        rom[169][23] = -8'd9;
        rom[169][24] = -8'd23;
        rom[169][25] = -8'd21;
        rom[169][26] = 8'd9;
        rom[169][27] = -8'd14;
        rom[169][28] = -8'd9;
        rom[169][29] = 8'd8;
        rom[169][30] = -8'd2;
        rom[169][31] = 8'd5;
        rom[169][32] = -8'd25;
        rom[169][33] = 8'd12;
        rom[169][34] = -8'd19;
        rom[169][35] = 8'd32;
        rom[169][36] = 8'd1;
        rom[169][37] = -8'd20;
        rom[169][38] = 8'd28;
        rom[169][39] = 8'd25;
        rom[169][40] = 8'd28;
        rom[169][41] = -8'd1;
        rom[169][42] = 8'd0;
        rom[169][43] = 8'd7;
        rom[169][44] = -8'd27;
        rom[169][45] = -8'd24;
        rom[169][46] = -8'd32;
        rom[169][47] = -8'd35;
        rom[169][48] = -8'd7;
        rom[169][49] = -8'd7;
        rom[169][50] = 8'd3;
        rom[169][51] = 8'd14;
        rom[169][52] = -8'd12;
        rom[169][53] = 8'd44;
        rom[169][54] = -8'd7;
        rom[169][55] = 8'd39;
        rom[169][56] = 8'd24;
        rom[169][57] = 8'd6;
        rom[169][58] = 8'd3;
        rom[169][59] = -8'd21;
        rom[169][60] = 8'd13;
        rom[169][61] = -8'd7;
        rom[169][62] = -8'd39;
        rom[169][63] = -8'd4;
        rom[170][0] = -8'd68;
        rom[170][1] = 8'd10;
        rom[170][2] = 8'd16;
        rom[170][3] = -8'd39;
        rom[170][4] = -8'd32;
        rom[170][5] = -8'd36;
        rom[170][6] = 8'd1;
        rom[170][7] = 8'd7;
        rom[170][8] = 8'd21;
        rom[170][9] = -8'd10;
        rom[170][10] = -8'd10;
        rom[170][11] = 8'd1;
        rom[170][12] = -8'd29;
        rom[170][13] = 8'd17;
        rom[170][14] = -8'd22;
        rom[170][15] = -8'd39;
        rom[170][16] = 8'd6;
        rom[170][17] = -8'd6;
        rom[170][18] = 8'd16;
        rom[170][19] = -8'd26;
        rom[170][20] = -8'd1;
        rom[170][21] = 8'd3;
        rom[170][22] = -8'd22;
        rom[170][23] = -8'd8;
        rom[170][24] = -8'd58;
        rom[170][25] = -8'd28;
        rom[170][26] = -8'd23;
        rom[170][27] = -8'd44;
        rom[170][28] = -8'd62;
        rom[170][29] = -8'd5;
        rom[170][30] = -8'd16;
        rom[170][31] = 8'd2;
        rom[170][32] = -8'd2;
        rom[170][33] = 8'd16;
        rom[170][34] = 8'd19;
        rom[170][35] = -8'd38;
        rom[170][36] = -8'd45;
        rom[170][37] = 8'd14;
        rom[170][38] = 8'd8;
        rom[170][39] = 8'd43;
        rom[170][40] = 8'd20;
        rom[170][41] = 8'd0;
        rom[170][42] = -8'd34;
        rom[170][43] = 8'd9;
        rom[170][44] = -8'd88;
        rom[170][45] = 8'd2;
        rom[170][46] = 8'd18;
        rom[170][47] = -8'd18;
        rom[170][48] = -8'd42;
        rom[170][49] = -8'd19;
        rom[170][50] = -8'd18;
        rom[170][51] = -8'd73;
        rom[170][52] = 8'd9;
        rom[170][53] = -8'd14;
        rom[170][54] = -8'd14;
        rom[170][55] = -8'd11;
        rom[170][56] = 8'd7;
        rom[170][57] = -8'd2;
        rom[170][58] = 8'd15;
        rom[170][59] = -8'd22;
        rom[170][60] = -8'd8;
        rom[170][61] = 8'd36;
        rom[170][62] = -8'd15;
        rom[170][63] = -8'd2;
        rom[171][0] = -8'd8;
        rom[171][1] = 8'd33;
        rom[171][2] = 8'd17;
        rom[171][3] = -8'd11;
        rom[171][4] = 8'd21;
        rom[171][5] = -8'd12;
        rom[171][6] = -8'd16;
        rom[171][7] = -8'd38;
        rom[171][8] = 8'd14;
        rom[171][9] = -8'd6;
        rom[171][10] = -8'd35;
        rom[171][11] = 8'd15;
        rom[171][12] = -8'd33;
        rom[171][13] = -8'd24;
        rom[171][14] = -8'd12;
        rom[171][15] = 8'd2;
        rom[171][16] = -8'd70;
        rom[171][17] = -8'd17;
        rom[171][18] = -8'd16;
        rom[171][19] = -8'd1;
        rom[171][20] = -8'd8;
        rom[171][21] = 8'd6;
        rom[171][22] = 8'd16;
        rom[171][23] = -8'd31;
        rom[171][24] = 8'd11;
        rom[171][25] = 8'd18;
        rom[171][26] = -8'd3;
        rom[171][27] = -8'd44;
        rom[171][28] = -8'd45;
        rom[171][29] = 8'd21;
        rom[171][30] = 8'd8;
        rom[171][31] = 8'd17;
        rom[171][32] = -8'd11;
        rom[171][33] = -8'd96;
        rom[171][34] = 8'd3;
        rom[171][35] = -8'd19;
        rom[171][36] = -8'd8;
        rom[171][37] = -8'd12;
        rom[171][38] = -8'd1;
        rom[171][39] = -8'd4;
        rom[171][40] = -8'd25;
        rom[171][41] = -8'd7;
        rom[171][42] = -8'd16;
        rom[171][43] = -8'd27;
        rom[171][44] = -8'd49;
        rom[171][45] = 8'd31;
        rom[171][46] = 8'd9;
        rom[171][47] = -8'd2;
        rom[171][48] = -8'd17;
        rom[171][49] = -8'd31;
        rom[171][50] = -8'd3;
        rom[171][51] = 8'd28;
        rom[171][52] = -8'd4;
        rom[171][53] = 8'd2;
        rom[171][54] = 8'd40;
        rom[171][55] = -8'd1;
        rom[171][56] = 8'd0;
        rom[171][57] = 8'd61;
        rom[171][58] = -8'd12;
        rom[171][59] = -8'd12;
        rom[171][60] = 8'd8;
        rom[171][61] = 8'd14;
        rom[171][62] = -8'd9;
        rom[171][63] = 8'd9;
        rom[172][0] = -8'd36;
        rom[172][1] = -8'd10;
        rom[172][2] = 8'd1;
        rom[172][3] = -8'd56;
        rom[172][4] = -8'd15;
        rom[172][5] = -8'd26;
        rom[172][6] = -8'd2;
        rom[172][7] = -8'd49;
        rom[172][8] = 8'd1;
        rom[172][9] = 8'd12;
        rom[172][10] = -8'd52;
        rom[172][11] = -8'd52;
        rom[172][12] = 8'd30;
        rom[172][13] = -8'd39;
        rom[172][14] = 8'd7;
        rom[172][15] = -8'd18;
        rom[172][16] = -8'd53;
        rom[172][17] = 8'd20;
        rom[172][18] = -8'd31;
        rom[172][19] = -8'd34;
        rom[172][20] = -8'd3;
        rom[172][21] = 8'd3;
        rom[172][22] = -8'd30;
        rom[172][23] = -8'd3;
        rom[172][24] = 8'd0;
        rom[172][25] = 8'd23;
        rom[172][26] = 8'd21;
        rom[172][27] = -8'd36;
        rom[172][28] = -8'd27;
        rom[172][29] = 8'd13;
        rom[172][30] = -8'd106;
        rom[172][31] = 8'd0;
        rom[172][32] = -8'd15;
        rom[172][33] = -8'd30;
        rom[172][34] = -8'd45;
        rom[172][35] = -8'd3;
        rom[172][36] = 8'd28;
        rom[172][37] = -8'd16;
        rom[172][38] = -8'd32;
        rom[172][39] = 8'd5;
        rom[172][40] = -8'd44;
        rom[172][41] = -8'd9;
        rom[172][42] = -8'd55;
        rom[172][43] = -8'd11;
        rom[172][44] = -8'd5;
        rom[172][45] = 8'd46;
        rom[172][46] = -8'd23;
        rom[172][47] = -8'd7;
        rom[172][48] = -8'd7;
        rom[172][49] = -8'd1;
        rom[172][50] = 8'd26;
        rom[172][51] = -8'd15;
        rom[172][52] = -8'd4;
        rom[172][53] = 8'd2;
        rom[172][54] = -8'd2;
        rom[172][55] = -8'd8;
        rom[172][56] = 8'd7;
        rom[172][57] = -8'd18;
        rom[172][58] = 8'd1;
        rom[172][59] = -8'd78;
        rom[172][60] = -8'd12;
        rom[172][61] = -8'd12;
        rom[172][62] = -8'd32;
        rom[172][63] = 8'd20;
        rom[173][0] = 8'd12;
        rom[173][1] = -8'd127;
        rom[173][2] = -8'd29;
        rom[173][3] = 8'd2;
        rom[173][4] = 8'd7;
        rom[173][5] = 8'd19;
        rom[173][6] = 8'd29;
        rom[173][7] = 8'd15;
        rom[173][8] = -8'd34;
        rom[173][9] = 8'd15;
        rom[173][10] = 8'd19;
        rom[173][11] = -8'd26;
        rom[173][12] = 8'd8;
        rom[173][13] = 8'd68;
        rom[173][14] = 8'd18;
        rom[173][15] = 8'd21;
        rom[173][16] = 8'd26;
        rom[173][17] = 8'd22;
        rom[173][18] = -8'd82;
        rom[173][19] = -8'd22;
        rom[173][20] = -8'd4;
        rom[173][21] = 8'd3;
        rom[173][22] = -8'd23;
        rom[173][23] = 8'd26;
        rom[173][24] = -8'd23;
        rom[173][25] = -8'd22;
        rom[173][26] = -8'd2;
        rom[173][27] = -8'd50;
        rom[173][28] = 8'd28;
        rom[173][29] = 8'd41;
        rom[173][30] = -8'd14;
        rom[173][31] = -8'd18;
        rom[173][32] = 8'd51;
        rom[173][33] = -8'd30;
        rom[173][34] = -8'd21;
        rom[173][35] = -8'd84;
        rom[173][36] = -8'd21;
        rom[173][37] = -8'd15;
        rom[173][38] = -8'd16;
        rom[173][39] = 8'd15;
        rom[173][40] = -8'd2;
        rom[173][41] = -8'd9;
        rom[173][42] = 8'd5;
        rom[173][43] = -8'd15;
        rom[173][44] = 8'd34;
        rom[173][45] = 8'd11;
        rom[173][46] = 8'd7;
        rom[173][47] = -8'd62;
        rom[173][48] = -8'd51;
        rom[173][49] = -8'd41;
        rom[173][50] = -8'd1;
        rom[173][51] = -8'd27;
        rom[173][52] = -8'd37;
        rom[173][53] = 8'd13;
        rom[173][54] = -8'd23;
        rom[173][55] = -8'd55;
        rom[173][56] = -8'd24;
        rom[173][57] = -8'd20;
        rom[173][58] = -8'd63;
        rom[173][59] = -8'd55;
        rom[173][60] = 8'd5;
        rom[173][61] = 8'd32;
        rom[173][62] = 8'd16;
        rom[173][63] = -8'd12;
        rom[174][0] = -8'd20;
        rom[174][1] = -8'd5;
        rom[174][2] = -8'd4;
        rom[174][3] = 8'd69;
        rom[174][4] = -8'd17;
        rom[174][5] = -8'd1;
        rom[174][6] = -8'd30;
        rom[174][7] = 8'd15;
        rom[174][8] = 8'd10;
        rom[174][9] = 8'd3;
        rom[174][10] = -8'd58;
        rom[174][11] = -8'd16;
        rom[174][12] = 8'd7;
        rom[174][13] = 8'd23;
        rom[174][14] = 8'd7;
        rom[174][15] = -8'd8;
        rom[174][16] = -8'd7;
        rom[174][17] = 8'd1;
        rom[174][18] = 8'd4;
        rom[174][19] = 8'd6;
        rom[174][20] = -8'd5;
        rom[174][21] = -8'd45;
        rom[174][22] = -8'd5;
        rom[174][23] = 8'd3;
        rom[174][24] = -8'd51;
        rom[174][25] = -8'd42;
        rom[174][26] = 8'd8;
        rom[174][27] = -8'd36;
        rom[174][28] = -8'd15;
        rom[174][29] = -8'd12;
        rom[174][30] = -8'd10;
        rom[174][31] = 8'd8;
        rom[174][32] = 8'd22;
        rom[174][33] = -8'd32;
        rom[174][34] = -8'd3;
        rom[174][35] = 8'd13;
        rom[174][36] = -8'd29;
        rom[174][37] = -8'd35;
        rom[174][38] = -8'd23;
        rom[174][39] = -8'd12;
        rom[174][40] = 8'd22;
        rom[174][41] = 8'd9;
        rom[174][42] = -8'd1;
        rom[174][43] = 8'd17;
        rom[174][44] = -8'd22;
        rom[174][45] = 8'd19;
        rom[174][46] = -8'd5;
        rom[174][47] = 8'd36;
        rom[174][48] = -8'd4;
        rom[174][49] = -8'd20;
        rom[174][50] = 8'd10;
        rom[174][51] = -8'd22;
        rom[174][52] = 8'd19;
        rom[174][53] = 8'd4;
        rom[174][54] = 8'd13;
        rom[174][55] = -8'd8;
        rom[174][56] = -8'd12;
        rom[174][57] = 8'd9;
        rom[174][58] = 8'd8;
        rom[174][59] = -8'd8;
        rom[174][60] = -8'd46;
        rom[174][61] = -8'd39;
        rom[174][62] = -8'd66;
        rom[174][63] = -8'd49;
        rom[175][0] = -8'd29;
        rom[175][1] = -8'd15;
        rom[175][2] = -8'd102;
        rom[175][3] = 8'd8;
        rom[175][4] = -8'd12;
        rom[175][5] = 8'd4;
        rom[175][6] = -8'd10;
        rom[175][7] = -8'd1;
        rom[175][8] = -8'd39;
        rom[175][9] = -8'd41;
        rom[175][10] = 8'd42;
        rom[175][11] = 8'd27;
        rom[175][12] = 8'd0;
        rom[175][13] = -8'd47;
        rom[175][14] = -8'd18;
        rom[175][15] = -8'd15;
        rom[175][16] = 8'd38;
        rom[175][17] = 8'd31;
        rom[175][18] = -8'd28;
        rom[175][19] = 8'd18;
        rom[175][20] = -8'd3;
        rom[175][21] = 8'd3;
        rom[175][22] = 8'd24;
        rom[175][23] = -8'd42;
        rom[175][24] = -8'd12;
        rom[175][25] = 8'd37;
        rom[175][26] = 8'd2;
        rom[175][27] = 8'd42;
        rom[175][28] = -8'd28;
        rom[175][29] = 8'd10;
        rom[175][30] = 8'd8;
        rom[175][31] = 8'd12;
        rom[175][32] = -8'd11;
        rom[175][33] = -8'd5;
        rom[175][34] = 8'd15;
        rom[175][35] = 8'd54;
        rom[175][36] = -8'd17;
        rom[175][37] = 8'd35;
        rom[175][38] = -8'd6;
        rom[175][39] = 8'd41;
        rom[175][40] = 8'd33;
        rom[175][41] = 8'd51;
        rom[175][42] = 8'd52;
        rom[175][43] = 8'd12;
        rom[175][44] = 8'd37;
        rom[175][45] = 8'd19;
        rom[175][46] = 8'd41;
        rom[175][47] = 8'd16;
        rom[175][48] = -8'd72;
        rom[175][49] = -8'd12;
        rom[175][50] = -8'd2;
        rom[175][51] = -8'd25;
        rom[175][52] = -8'd5;
        rom[175][53] = -8'd20;
        rom[175][54] = 8'd15;
        rom[175][55] = -8'd10;
        rom[175][56] = -8'd9;
        rom[175][57] = -8'd34;
        rom[175][58] = -8'd27;
        rom[175][59] = -8'd16;
        rom[175][60] = -8'd26;
        rom[175][61] = -8'd71;
        rom[175][62] = -8'd13;
        rom[175][63] = 8'd5;
        rom[176][0] = -8'd51;
        rom[176][1] = 8'd3;
        rom[176][2] = -8'd36;
        rom[176][3] = 8'd49;
        rom[176][4] = -8'd2;
        rom[176][5] = 8'd25;
        rom[176][6] = -8'd83;
        rom[176][7] = -8'd20;
        rom[176][8] = -8'd5;
        rom[176][9] = -8'd16;
        rom[176][10] = -8'd34;
        rom[176][11] = 8'd18;
        rom[176][12] = 8'd14;
        rom[176][13] = -8'd9;
        rom[176][14] = -8'd1;
        rom[176][15] = 8'd46;
        rom[176][16] = 8'd34;
        rom[176][17] = -8'd49;
        rom[176][18] = -8'd45;
        rom[176][19] = -8'd22;
        rom[176][20] = -8'd9;
        rom[176][21] = -8'd2;
        rom[176][22] = -8'd80;
        rom[176][23] = -8'd59;
        rom[176][24] = -8'd10;
        rom[176][25] = -8'd14;
        rom[176][26] = -8'd29;
        rom[176][27] = -8'd36;
        rom[176][28] = 8'd11;
        rom[176][29] = -8'd55;
        rom[176][30] = 8'd4;
        rom[176][31] = 8'd9;
        rom[176][32] = -8'd2;
        rom[176][33] = -8'd22;
        rom[176][34] = 8'd14;
        rom[176][35] = -8'd32;
        rom[176][36] = -8'd23;
        rom[176][37] = -8'd28;
        rom[176][38] = -8'd58;
        rom[176][39] = 8'd7;
        rom[176][40] = 8'd23;
        rom[176][41] = -8'd34;
        rom[176][42] = -8'd3;
        rom[176][43] = 8'd29;
        rom[176][44] = 8'd5;
        rom[176][45] = -8'd29;
        rom[176][46] = 8'd2;
        rom[176][47] = -8'd2;
        rom[176][48] = -8'd88;
        rom[176][49] = -8'd11;
        rom[176][50] = -8'd10;
        rom[176][51] = -8'd66;
        rom[176][52] = 8'd28;
        rom[176][53] = -8'd53;
        rom[176][54] = -8'd5;
        rom[176][55] = -8'd3;
        rom[176][56] = 8'd4;
        rom[176][57] = -8'd7;
        rom[176][58] = -8'd20;
        rom[176][59] = 8'd2;
        rom[176][60] = -8'd27;
        rom[176][61] = -8'd47;
        rom[176][62] = -8'd19;
        rom[176][63] = -8'd46;
        rom[177][0] = -8'd40;
        rom[177][1] = 8'd8;
        rom[177][2] = 8'd7;
        rom[177][3] = 8'd6;
        rom[177][4] = -8'd3;
        rom[177][5] = -8'd5;
        rom[177][6] = -8'd20;
        rom[177][7] = -8'd57;
        rom[177][8] = 8'd17;
        rom[177][9] = 8'd10;
        rom[177][10] = -8'd33;
        rom[177][11] = 8'd11;
        rom[177][12] = 8'd27;
        rom[177][13] = -8'd8;
        rom[177][14] = -8'd25;
        rom[177][15] = -8'd15;
        rom[177][16] = 8'd26;
        rom[177][17] = -8'd13;
        rom[177][18] = -8'd31;
        rom[177][19] = 8'd0;
        rom[177][20] = 8'd0;
        rom[177][21] = -8'd9;
        rom[177][22] = 8'd26;
        rom[177][23] = -8'd26;
        rom[177][24] = 8'd37;
        rom[177][25] = -8'd4;
        rom[177][26] = -8'd21;
        rom[177][27] = 8'd49;
        rom[177][28] = 8'd45;
        rom[177][29] = 8'd19;
        rom[177][30] = 8'd15;
        rom[177][31] = 8'd21;
        rom[177][32] = -8'd7;
        rom[177][33] = -8'd18;
        rom[177][34] = 8'd17;
        rom[177][35] = 8'd29;
        rom[177][36] = -8'd27;
        rom[177][37] = 8'd15;
        rom[177][38] = -8'd30;
        rom[177][39] = -8'd17;
        rom[177][40] = -8'd15;
        rom[177][41] = -8'd5;
        rom[177][42] = -8'd62;
        rom[177][43] = -8'd3;
        rom[177][44] = -8'd1;
        rom[177][45] = -8'd4;
        rom[177][46] = -8'd5;
        rom[177][47] = 8'd24;
        rom[177][48] = 8'd10;
        rom[177][49] = -8'd2;
        rom[177][50] = 8'd9;
        rom[177][51] = -8'd4;
        rom[177][52] = -8'd51;
        rom[177][53] = -8'd2;
        rom[177][54] = 8'd18;
        rom[177][55] = 8'd18;
        rom[177][56] = -8'd31;
        rom[177][57] = -8'd26;
        rom[177][58] = -8'd22;
        rom[177][59] = 8'd19;
        rom[177][60] = 8'd43;
        rom[177][61] = -8'd19;
        rom[177][62] = 8'd1;
        rom[177][63] = 8'd10;
        rom[178][0] = 8'd23;
        rom[178][1] = -8'd1;
        rom[178][2] = 8'd0;
        rom[178][3] = 8'd13;
        rom[178][4] = -8'd26;
        rom[178][5] = 8'd29;
        rom[178][6] = -8'd9;
        rom[178][7] = -8'd6;
        rom[178][8] = -8'd26;
        rom[178][9] = -8'd16;
        rom[178][10] = -8'd41;
        rom[178][11] = -8'd16;
        rom[178][12] = 8'd27;
        rom[178][13] = 8'd10;
        rom[178][14] = 8'd25;
        rom[178][15] = -8'd52;
        rom[178][16] = -8'd19;
        rom[178][17] = 8'd20;
        rom[178][18] = -8'd3;
        rom[178][19] = -8'd6;
        rom[178][20] = 8'd0;
        rom[178][21] = -8'd47;
        rom[178][22] = 8'd21;
        rom[178][23] = 8'd5;
        rom[178][24] = -8'd16;
        rom[178][25] = -8'd59;
        rom[178][26] = -8'd17;
        rom[178][27] = 8'd42;
        rom[178][28] = -8'd41;
        rom[178][29] = -8'd14;
        rom[178][30] = -8'd9;
        rom[178][31] = -8'd21;
        rom[178][32] = 8'd11;
        rom[178][33] = 8'd32;
        rom[178][34] = -8'd32;
        rom[178][35] = -8'd5;
        rom[178][36] = 8'd8;
        rom[178][37] = 8'd13;
        rom[178][38] = 8'd3;
        rom[178][39] = -8'd23;
        rom[178][40] = -8'd4;
        rom[178][41] = 8'd45;
        rom[178][42] = 8'd30;
        rom[178][43] = -8'd54;
        rom[178][44] = -8'd7;
        rom[178][45] = -8'd31;
        rom[178][46] = -8'd25;
        rom[178][47] = 8'd7;
        rom[178][48] = 8'd11;
        rom[178][49] = 8'd6;
        rom[178][50] = 8'd27;
        rom[178][51] = -8'd50;
        rom[178][52] = 8'd18;
        rom[178][53] = -8'd67;
        rom[178][54] = -8'd24;
        rom[178][55] = 8'd21;
        rom[178][56] = -8'd2;
        rom[178][57] = 8'd1;
        rom[178][58] = -8'd8;
        rom[178][59] = 8'd2;
        rom[178][60] = -8'd42;
        rom[178][61] = -8'd10;
        rom[178][62] = -8'd33;
        rom[178][63] = -8'd10;
        rom[179][0] = 8'd30;
        rom[179][1] = 8'd11;
        rom[179][2] = 8'd26;
        rom[179][3] = 8'd1;
        rom[179][4] = 8'd15;
        rom[179][5] = -8'd41;
        rom[179][6] = -8'd9;
        rom[179][7] = -8'd5;
        rom[179][8] = 8'd15;
        rom[179][9] = 8'd33;
        rom[179][10] = 8'd24;
        rom[179][11] = 8'd18;
        rom[179][12] = -8'd21;
        rom[179][13] = -8'd13;
        rom[179][14] = 8'd15;
        rom[179][15] = 8'd36;
        rom[179][16] = -8'd26;
        rom[179][17] = -8'd7;
        rom[179][18] = -8'd19;
        rom[179][19] = 8'd14;
        rom[179][20] = 8'd4;
        rom[179][21] = -8'd24;
        rom[179][22] = -8'd24;
        rom[179][23] = -8'd6;
        rom[179][24] = -8'd49;
        rom[179][25] = -8'd23;
        rom[179][26] = 8'd1;
        rom[179][27] = 8'd28;
        rom[179][28] = -8'd11;
        rom[179][29] = -8'd1;
        rom[179][30] = 8'd15;
        rom[179][31] = -8'd5;
        rom[179][32] = 8'd10;
        rom[179][33] = 8'd57;
        rom[179][34] = -8'd24;
        rom[179][35] = 8'd43;
        rom[179][36] = 8'd12;
        rom[179][37] = 8'd42;
        rom[179][38] = -8'd11;
        rom[179][39] = 8'd12;
        rom[179][40] = -8'd40;
        rom[179][41] = -8'd19;
        rom[179][42] = 8'd26;
        rom[179][43] = -8'd39;
        rom[179][44] = 8'd2;
        rom[179][45] = 8'd14;
        rom[179][46] = 8'd63;
        rom[179][47] = -8'd19;
        rom[179][48] = -8'd4;
        rom[179][49] = -8'd9;
        rom[179][50] = 8'd30;
        rom[179][51] = -8'd18;
        rom[179][52] = -8'd64;
        rom[179][53] = -8'd30;
        rom[179][54] = -8'd2;
        rom[179][55] = 8'd2;
        rom[179][56] = -8'd15;
        rom[179][57] = 8'd0;
        rom[179][58] = -8'd11;
        rom[179][59] = -8'd43;
        rom[179][60] = 8'd7;
        rom[179][61] = 8'd15;
        rom[179][62] = 8'd6;
        rom[179][63] = -8'd18;
        rom[180][0] = -8'd24;
        rom[180][1] = -8'd6;
        rom[180][2] = 8'd12;
        rom[180][3] = -8'd3;
        rom[180][4] = 8'd5;
        rom[180][5] = -8'd33;
        rom[180][6] = -8'd43;
        rom[180][7] = -8'd12;
        rom[180][8] = 8'd12;
        rom[180][9] = -8'd5;
        rom[180][10] = -8'd13;
        rom[180][11] = 8'd16;
        rom[180][12] = -8'd75;
        rom[180][13] = 8'd49;
        rom[180][14] = 8'd13;
        rom[180][15] = -8'd5;
        rom[180][16] = 8'd2;
        rom[180][17] = 8'd6;
        rom[180][18] = 8'd9;
        rom[180][19] = -8'd46;
        rom[180][20] = 8'd0;
        rom[180][21] = -8'd6;
        rom[180][22] = 8'd19;
        rom[180][23] = -8'd12;
        rom[180][24] = -8'd8;
        rom[180][25] = 8'd6;
        rom[180][26] = -8'd8;
        rom[180][27] = -8'd36;
        rom[180][28] = -8'd4;
        rom[180][29] = -8'd6;
        rom[180][30] = -8'd14;
        rom[180][31] = 8'd10;
        rom[180][32] = -8'd4;
        rom[180][33] = -8'd3;
        rom[180][34] = 8'd27;
        rom[180][35] = -8'd1;
        rom[180][36] = -8'd8;
        rom[180][37] = -8'd8;
        rom[180][38] = 8'd25;
        rom[180][39] = 8'd3;
        rom[180][40] = -8'd19;
        rom[180][41] = 8'd23;
        rom[180][42] = 8'd68;
        rom[180][43] = 8'd10;
        rom[180][44] = -8'd14;
        rom[180][45] = -8'd65;
        rom[180][46] = -8'd43;
        rom[180][47] = -8'd52;
        rom[180][48] = 8'd18;
        rom[180][49] = 8'd5;
        rom[180][50] = 8'd4;
        rom[180][51] = -8'd10;
        rom[180][52] = 8'd5;
        rom[180][53] = 8'd13;
        rom[180][54] = -8'd45;
        rom[180][55] = 8'd3;
        rom[180][56] = -8'd9;
        rom[180][57] = 8'd12;
        rom[180][58] = -8'd10;
        rom[180][59] = 8'd1;
        rom[180][60] = -8'd31;
        rom[180][61] = 8'd19;
        rom[180][62] = 8'd10;
        rom[180][63] = 8'd10;
        rom[181][0] = -8'd30;
        rom[181][1] = -8'd9;
        rom[181][2] = -8'd47;
        rom[181][3] = -8'd6;
        rom[181][4] = 8'd3;
        rom[181][5] = -8'd13;
        rom[181][6] = 8'd0;
        rom[181][7] = -8'd1;
        rom[181][8] = 8'd1;
        rom[181][9] = -8'd2;
        rom[181][10] = 8'd17;
        rom[181][11] = -8'd1;
        rom[181][12] = 8'd42;
        rom[181][13] = 8'd9;
        rom[181][14] = -8'd23;
        rom[181][15] = 8'd31;
        rom[181][16] = 8'd23;
        rom[181][17] = 8'd3;
        rom[181][18] = -8'd11;
        rom[181][19] = -8'd52;
        rom[181][20] = -8'd5;
        rom[181][21] = 8'd23;
        rom[181][22] = 8'd6;
        rom[181][23] = -8'd27;
        rom[181][24] = -8'd36;
        rom[181][25] = -8'd7;
        rom[181][26] = 8'd3;
        rom[181][27] = -8'd19;
        rom[181][28] = 8'd3;
        rom[181][29] = -8'd29;
        rom[181][30] = 8'd17;
        rom[181][31] = 8'd26;
        rom[181][32] = 8'd22;
        rom[181][33] = -8'd51;
        rom[181][34] = 8'd15;
        rom[181][35] = 8'd19;
        rom[181][36] = -8'd47;
        rom[181][37] = -8'd49;
        rom[181][38] = 8'd3;
        rom[181][39] = 8'd3;
        rom[181][40] = 8'd30;
        rom[181][41] = -8'd3;
        rom[181][42] = 8'd7;
        rom[181][43] = 8'd17;
        rom[181][44] = -8'd31;
        rom[181][45] = -8'd34;
        rom[181][46] = -8'd4;
        rom[181][47] = -8'd10;
        rom[181][48] = -8'd49;
        rom[181][49] = -8'd3;
        rom[181][50] = -8'd72;
        rom[181][51] = -8'd8;
        rom[181][52] = -8'd2;
        rom[181][53] = 8'd32;
        rom[181][54] = 8'd9;
        rom[181][55] = -8'd23;
        rom[181][56] = 8'd9;
        rom[181][57] = -8'd3;
        rom[181][58] = -8'd41;
        rom[181][59] = -8'd16;
        rom[181][60] = 8'd10;
        rom[181][61] = -8'd18;
        rom[181][62] = -8'd43;
        rom[181][63] = -8'd15;
        rom[182][0] = 8'd9;
        rom[182][1] = -8'd5;
        rom[182][2] = 8'd1;
        rom[182][3] = -8'd7;
        rom[182][4] = -8'd1;
        rom[182][5] = -8'd5;
        rom[182][6] = -8'd4;
        rom[182][7] = -8'd1;
        rom[182][8] = 8'd8;
        rom[182][9] = -8'd5;
        rom[182][10] = 8'd3;
        rom[182][11] = 8'd7;
        rom[182][12] = 8'd8;
        rom[182][13] = -8'd1;
        rom[182][14] = -8'd1;
        rom[182][15] = -8'd7;
        rom[182][16] = -8'd10;
        rom[182][17] = 8'd8;
        rom[182][18] = 8'd1;
        rom[182][19] = 8'd4;
        rom[182][20] = -8'd2;
        rom[182][21] = -8'd8;
        rom[182][22] = -8'd6;
        rom[182][23] = -8'd2;
        rom[182][24] = 8'd8;
        rom[182][25] = -8'd9;
        rom[182][26] = 8'd11;
        rom[182][27] = 8'd6;
        rom[182][28] = 8'd8;
        rom[182][29] = -8'd4;
        rom[182][30] = -8'd6;
        rom[182][31] = 8'd10;
        rom[182][32] = -8'd7;
        rom[182][33] = -8'd7;
        rom[182][34] = 8'd9;
        rom[182][35] = 8'd6;
        rom[182][36] = -8'd8;
        rom[182][37] = 8'd2;
        rom[182][38] = -8'd9;
        rom[182][39] = 8'd0;
        rom[182][40] = -8'd3;
        rom[182][41] = 8'd8;
        rom[182][42] = -8'd8;
        rom[182][43] = -8'd8;
        rom[182][44] = -8'd1;
        rom[182][45] = 8'd3;
        rom[182][46] = -8'd2;
        rom[182][47] = -8'd6;
        rom[182][48] = 8'd0;
        rom[182][49] = 8'd1;
        rom[182][50] = -8'd6;
        rom[182][51] = -8'd9;
        rom[182][52] = 8'd1;
        rom[182][53] = 8'd1;
        rom[182][54] = 8'd4;
        rom[182][55] = -8'd7;
        rom[182][56] = -8'd6;
        rom[182][57] = -8'd3;
        rom[182][58] = -8'd7;
        rom[182][59] = -8'd5;
        rom[182][60] = -8'd7;
        rom[182][61] = -8'd10;
        rom[182][62] = 8'd2;
        rom[182][63] = 8'd5;
        rom[183][0] = -8'd25;
        rom[183][1] = 8'd21;
        rom[183][2] = -8'd26;
        rom[183][3] = 8'd8;
        rom[183][4] = -8'd19;
        rom[183][5] = 8'd29;
        rom[183][6] = 8'd12;
        rom[183][7] = 8'd18;
        rom[183][8] = 8'd32;
        rom[183][9] = 8'd17;
        rom[183][10] = -8'd24;
        rom[183][11] = -8'd31;
        rom[183][12] = -8'd22;
        rom[183][13] = 8'd13;
        rom[183][14] = -8'd9;
        rom[183][15] = 8'd2;
        rom[183][16] = 8'd10;
        rom[183][17] = 8'd6;
        rom[183][18] = 8'd12;
        rom[183][19] = 8'd14;
        rom[183][20] = -8'd18;
        rom[183][21] = 8'd63;
        rom[183][22] = -8'd88;
        rom[183][23] = -8'd109;
        rom[183][24] = 8'd2;
        rom[183][25] = -8'd4;
        rom[183][26] = -8'd32;
        rom[183][27] = -8'd18;
        rom[183][28] = 8'd2;
        rom[183][29] = 8'd56;
        rom[183][30] = 8'd23;
        rom[183][31] = 8'd34;
        rom[183][32] = 8'd12;
        rom[183][33] = 8'd37;
        rom[183][34] = -8'd17;
        rom[183][35] = 8'd11;
        rom[183][36] = 8'd27;
        rom[183][37] = -8'd9;
        rom[183][38] = 8'd24;
        rom[183][39] = 8'd19;
        rom[183][40] = 8'd57;
        rom[183][41] = 8'd16;
        rom[183][42] = -8'd26;
        rom[183][43] = 8'd20;
        rom[183][44] = -8'd40;
        rom[183][45] = 8'd17;
        rom[183][46] = 8'd20;
        rom[183][47] = -8'd63;
        rom[183][48] = -8'd29;
        rom[183][49] = 8'd10;
        rom[183][50] = -8'd37;
        rom[183][51] = -8'd15;
        rom[183][52] = 8'd17;
        rom[183][53] = 8'd40;
        rom[183][54] = -8'd69;
        rom[183][55] = 8'd16;
        rom[183][56] = -8'd59;
        rom[183][57] = -8'd3;
        rom[183][58] = 8'd19;
        rom[183][59] = 8'd14;
        rom[183][60] = 8'd12;
        rom[183][61] = 8'd8;
        rom[183][62] = -8'd3;
        rom[183][63] = 8'd6;
        rom[184][0] = -8'd48;
        rom[184][1] = -8'd10;
        rom[184][2] = -8'd7;
        rom[184][3] = -8'd15;
        rom[184][4] = 8'd2;
        rom[184][5] = -8'd79;
        rom[184][6] = -8'd70;
        rom[184][7] = -8'd49;
        rom[184][8] = -8'd23;
        rom[184][9] = -8'd35;
        rom[184][10] = 8'd18;
        rom[184][11] = -8'd27;
        rom[184][12] = 8'd23;
        rom[184][13] = -8'd55;
        rom[184][14] = 8'd18;
        rom[184][15] = -8'd20;
        rom[184][16] = 8'd20;
        rom[184][17] = 8'd36;
        rom[184][18] = -8'd42;
        rom[184][19] = -8'd47;
        rom[184][20] = -8'd8;
        rom[184][21] = -8'd25;
        rom[184][22] = 8'd41;
        rom[184][23] = -8'd58;
        rom[184][24] = 8'd3;
        rom[184][25] = -8'd4;
        rom[184][26] = 8'd2;
        rom[184][27] = -8'd9;
        rom[184][28] = -8'd11;
        rom[184][29] = 8'd18;
        rom[184][30] = -8'd80;
        rom[184][31] = 8'd5;
        rom[184][32] = -8'd35;
        rom[184][33] = -8'd66;
        rom[184][34] = -8'd4;
        rom[184][35] = 8'd31;
        rom[184][36] = 8'd17;
        rom[184][37] = 8'd14;
        rom[184][38] = -8'd34;
        rom[184][39] = -8'd34;
        rom[184][40] = 8'd13;
        rom[184][41] = 8'd3;
        rom[184][42] = 8'd6;
        rom[184][43] = 8'd28;
        rom[184][44] = -8'd23;
        rom[184][45] = -8'd50;
        rom[184][46] = 8'd20;
        rom[184][47] = -8'd39;
        rom[184][48] = -8'd57;
        rom[184][49] = -8'd8;
        rom[184][50] = 8'd30;
        rom[184][51] = -8'd12;
        rom[184][52] = 8'd9;
        rom[184][53] = 8'd26;
        rom[184][54] = -8'd30;
        rom[184][55] = 8'd10;
        rom[184][56] = -8'd15;
        rom[184][57] = -8'd16;
        rom[184][58] = -8'd32;
        rom[184][59] = -8'd45;
        rom[184][60] = -8'd9;
        rom[184][61] = 8'd34;
        rom[184][62] = -8'd19;
        rom[184][63] = 8'd0;
        rom[185][0] = -8'd35;
        rom[185][1] = -8'd40;
        rom[185][2] = 8'd1;
        rom[185][3] = -8'd7;
        rom[185][4] = 8'd33;
        rom[185][5] = 8'd35;
        rom[185][6] = 8'd5;
        rom[185][7] = 8'd1;
        rom[185][8] = -8'd16;
        rom[185][9] = 8'd25;
        rom[185][10] = -8'd37;
        rom[185][11] = -8'd30;
        rom[185][12] = -8'd10;
        rom[185][13] = 8'd4;
        rom[185][14] = 8'd18;
        rom[185][15] = -8'd13;
        rom[185][16] = -8'd22;
        rom[185][17] = 8'd11;
        rom[185][18] = -8'd24;
        rom[185][19] = 8'd14;
        rom[185][20] = -8'd7;
        rom[185][21] = 8'd7;
        rom[185][22] = -8'd7;
        rom[185][23] = -8'd8;
        rom[185][24] = 8'd12;
        rom[185][25] = 8'd9;
        rom[185][26] = -8'd3;
        rom[185][27] = -8'd26;
        rom[185][28] = 8'd32;
        rom[185][29] = 8'd28;
        rom[185][30] = -8'd1;
        rom[185][31] = 8'd5;
        rom[185][32] = 8'd8;
        rom[185][33] = 8'd14;
        rom[185][34] = 8'd24;
        rom[185][35] = 8'd1;
        rom[185][36] = 8'd47;
        rom[185][37] = -8'd37;
        rom[185][38] = -8'd3;
        rom[185][39] = 8'd11;
        rom[185][40] = -8'd20;
        rom[185][41] = 8'd17;
        rom[185][42] = 8'd10;
        rom[185][43] = -8'd77;
        rom[185][44] = 8'd43;
        rom[185][45] = 8'd15;
        rom[185][46] = 8'd1;
        rom[185][47] = 8'd8;
        rom[185][48] = 8'd21;
        rom[185][49] = -8'd24;
        rom[185][50] = -8'd16;
        rom[185][51] = -8'd8;
        rom[185][52] = 8'd16;
        rom[185][53] = -8'd12;
        rom[185][54] = 8'd43;
        rom[185][55] = -8'd5;
        rom[185][56] = 8'd6;
        rom[185][57] = -8'd2;
        rom[185][58] = -8'd22;
        rom[185][59] = -8'd6;
        rom[185][60] = 8'd21;
        rom[185][61] = 8'd15;
        rom[185][62] = -8'd44;
        rom[185][63] = 8'd14;
        rom[186][0] = 8'd10;
        rom[186][1] = -8'd37;
        rom[186][2] = -8'd11;
        rom[186][3] = 8'd39;
        rom[186][4] = -8'd29;
        rom[186][5] = 8'd0;
        rom[186][6] = 8'd14;
        rom[186][7] = 8'd17;
        rom[186][8] = -8'd45;
        rom[186][9] = 8'd2;
        rom[186][10] = -8'd11;
        rom[186][11] = -8'd6;
        rom[186][12] = -8'd52;
        rom[186][13] = -8'd53;
        rom[186][14] = 8'd42;
        rom[186][15] = 8'd10;
        rom[186][16] = -8'd10;
        rom[186][17] = -8'd52;
        rom[186][18] = -8'd36;
        rom[186][19] = 8'd9;
        rom[186][20] = -8'd10;
        rom[186][21] = 8'd68;
        rom[186][22] = 8'd0;
        rom[186][23] = -8'd55;
        rom[186][24] = -8'd32;
        rom[186][25] = 8'd6;
        rom[186][26] = 8'd29;
        rom[186][27] = -8'd14;
        rom[186][28] = -8'd36;
        rom[186][29] = -8'd40;
        rom[186][30] = 8'd33;
        rom[186][31] = -8'd42;
        rom[186][32] = -8'd28;
        rom[186][33] = -8'd35;
        rom[186][34] = 8'd8;
        rom[186][35] = -8'd18;
        rom[186][36] = 8'd1;
        rom[186][37] = 8'd7;
        rom[186][38] = 8'd37;
        rom[186][39] = -8'd1;
        rom[186][40] = 8'd16;
        rom[186][41] = -8'd3;
        rom[186][42] = -8'd14;
        rom[186][43] = -8'd5;
        rom[186][44] = 8'd1;
        rom[186][45] = -8'd36;
        rom[186][46] = -8'd2;
        rom[186][47] = -8'd47;
        rom[186][48] = 8'd62;
        rom[186][49] = 8'd3;
        rom[186][50] = 8'd14;
        rom[186][51] = 8'd21;
        rom[186][52] = -8'd5;
        rom[186][53] = 8'd15;
        rom[186][54] = 8'd3;
        rom[186][55] = 8'd15;
        rom[186][56] = 8'd39;
        rom[186][57] = -8'd58;
        rom[186][58] = 8'd44;
        rom[186][59] = 8'd65;
        rom[186][60] = 8'd28;
        rom[186][61] = 8'd5;
        rom[186][62] = -8'd34;
        rom[186][63] = -8'd5;
        rom[187][0] = -8'd11;
        rom[187][1] = -8'd54;
        rom[187][2] = -8'd4;
        rom[187][3] = 8'd7;
        rom[187][4] = -8'd6;
        rom[187][5] = 8'd10;
        rom[187][6] = -8'd127;
        rom[187][7] = -8'd9;
        rom[187][8] = 8'd20;
        rom[187][9] = 8'd6;
        rom[187][10] = -8'd26;
        rom[187][11] = -8'd19;
        rom[187][12] = 8'd5;
        rom[187][13] = -8'd33;
        rom[187][14] = 8'd15;
        rom[187][15] = -8'd9;
        rom[187][16] = 8'd5;
        rom[187][17] = -8'd25;
        rom[187][18] = -8'd48;
        rom[187][19] = -8'd7;
        rom[187][20] = -8'd1;
        rom[187][21] = 8'd26;
        rom[187][22] = -8'd6;
        rom[187][23] = -8'd15;
        rom[187][24] = 8'd5;
        rom[187][25] = 8'd7;
        rom[187][26] = -8'd21;
        rom[187][27] = -8'd39;
        rom[187][28] = 8'd20;
        rom[187][29] = -8'd4;
        rom[187][30] = -8'd49;
        rom[187][31] = -8'd20;
        rom[187][32] = -8'd46;
        rom[187][33] = -8'd62;
        rom[187][34] = 8'd14;
        rom[187][35] = -8'd13;
        rom[187][36] = -8'd6;
        rom[187][37] = -8'd16;
        rom[187][38] = 8'd9;
        rom[187][39] = -8'd10;
        rom[187][40] = -8'd1;
        rom[187][41] = -8'd8;
        rom[187][42] = -8'd6;
        rom[187][43] = 8'd14;
        rom[187][44] = -8'd38;
        rom[187][45] = 8'd30;
        rom[187][46] = 8'd16;
        rom[187][47] = 8'd15;
        rom[187][48] = 8'd22;
        rom[187][49] = 8'd17;
        rom[187][50] = 8'd25;
        rom[187][51] = -8'd11;
        rom[187][52] = -8'd18;
        rom[187][53] = -8'd27;
        rom[187][54] = 8'd19;
        rom[187][55] = 8'd4;
        rom[187][56] = -8'd98;
        rom[187][57] = 8'd4;
        rom[187][58] = 8'd14;
        rom[187][59] = -8'd43;
        rom[187][60] = -8'd33;
        rom[187][61] = 8'd28;
        rom[187][62] = 8'd2;
        rom[187][63] = 8'd9;
        rom[188][0] = -8'd22;
        rom[188][1] = 8'd27;
        rom[188][2] = -8'd19;
        rom[188][3] = -8'd39;
        rom[188][4] = -8'd9;
        rom[188][5] = -8'd44;
        rom[188][6] = -8'd14;
        rom[188][7] = 8'd26;
        rom[188][8] = 8'd11;
        rom[188][9] = -8'd22;
        rom[188][10] = -8'd22;
        rom[188][11] = -8'd29;
        rom[188][12] = 8'd25;
        rom[188][13] = -8'd5;
        rom[188][14] = 8'd16;
        rom[188][15] = 8'd19;
        rom[188][16] = -8'd34;
        rom[188][17] = -8'd6;
        rom[188][18] = -8'd13;
        rom[188][19] = -8'd4;
        rom[188][20] = -8'd9;
        rom[188][21] = -8'd58;
        rom[188][22] = 8'd11;
        rom[188][23] = 8'd5;
        rom[188][24] = -8'd24;
        rom[188][25] = -8'd19;
        rom[188][26] = -8'd13;
        rom[188][27] = 8'd51;
        rom[188][28] = 8'd3;
        rom[188][29] = -8'd11;
        rom[188][30] = 8'd22;
        rom[188][31] = -8'd32;
        rom[188][32] = 8'd30;
        rom[188][33] = 8'd38;
        rom[188][34] = -8'd39;
        rom[188][35] = 8'd18;
        rom[188][36] = -8'd8;
        rom[188][37] = 8'd21;
        rom[188][38] = 8'd4;
        rom[188][39] = 8'd4;
        rom[188][40] = -8'd6;
        rom[188][41] = 8'd1;
        rom[188][42] = 8'd0;
        rom[188][43] = 8'd31;
        rom[188][44] = 8'd40;
        rom[188][45] = 8'd28;
        rom[188][46] = -8'd36;
        rom[188][47] = -8'd82;
        rom[188][48] = -8'd16;
        rom[188][49] = 8'd46;
        rom[188][50] = 8'd3;
        rom[188][51] = -8'd30;
        rom[188][52] = 8'd45;
        rom[188][53] = -8'd19;
        rom[188][54] = -8'd22;
        rom[188][55] = -8'd3;
        rom[188][56] = -8'd6;
        rom[188][57] = 8'd69;
        rom[188][58] = 8'd38;
        rom[188][59] = -8'd15;
        rom[188][60] = -8'd46;
        rom[188][61] = -8'd1;
        rom[188][62] = -8'd26;
        rom[188][63] = -8'd4;
        rom[189][0] = -8'd14;
        rom[189][1] = 8'd0;
        rom[189][2] = 8'd17;
        rom[189][3] = -8'd23;
        rom[189][4] = -8'd4;
        rom[189][5] = -8'd21;
        rom[189][6] = 8'd33;
        rom[189][7] = -8'd8;
        rom[189][8] = -8'd16;
        rom[189][9] = 8'd17;
        rom[189][10] = -8'd50;
        rom[189][11] = 8'd12;
        rom[189][12] = 8'd9;
        rom[189][13] = -8'd26;
        rom[189][14] = 8'd8;
        rom[189][15] = 8'd4;
        rom[189][16] = 8'd1;
        rom[189][17] = 8'd16;
        rom[189][18] = 8'd10;
        rom[189][19] = 8'd0;
        rom[189][20] = -8'd4;
        rom[189][21] = 8'd20;
        rom[189][22] = 8'd33;
        rom[189][23] = -8'd47;
        rom[189][24] = 8'd18;
        rom[189][25] = -8'd21;
        rom[189][26] = -8'd64;
        rom[189][27] = 8'd0;
        rom[189][28] = -8'd11;
        rom[189][29] = 8'd27;
        rom[189][30] = -8'd70;
        rom[189][31] = -8'd16;
        rom[189][32] = -8'd12;
        rom[189][33] = 8'd23;
        rom[189][34] = -8'd2;
        rom[189][35] = 8'd36;
        rom[189][36] = 8'd11;
        rom[189][37] = 8'd18;
        rom[189][38] = -8'd42;
        rom[189][39] = 8'd1;
        rom[189][40] = -8'd43;
        rom[189][41] = 8'd12;
        rom[189][42] = -8'd36;
        rom[189][43] = -8'd52;
        rom[189][44] = 8'd18;
        rom[189][45] = 8'd20;
        rom[189][46] = -8'd9;
        rom[189][47] = 8'd26;
        rom[189][48] = -8'd20;
        rom[189][49] = 8'd22;
        rom[189][50] = 8'd24;
        rom[189][51] = -8'd8;
        rom[189][52] = -8'd23;
        rom[189][53] = -8'd16;
        rom[189][54] = -8'd31;
        rom[189][55] = 8'd21;
        rom[189][56] = -8'd2;
        rom[189][57] = -8'd18;
        rom[189][58] = -8'd30;
        rom[189][59] = -8'd87;
        rom[189][60] = 8'd58;
        rom[189][61] = -8'd79;
        rom[189][62] = -8'd6;
        rom[189][63] = 8'd30;
        rom[190][0] = 8'd9;
        rom[190][1] = -8'd20;
        rom[190][2] = 8'd8;
        rom[190][3] = -8'd57;
        rom[190][4] = -8'd33;
        rom[190][5] = -8'd31;
        rom[190][6] = -8'd51;
        rom[190][7] = 8'd15;
        rom[190][8] = -8'd33;
        rom[190][9] = 8'd12;
        rom[190][10] = -8'd36;
        rom[190][11] = 8'd13;
        rom[190][12] = 8'd41;
        rom[190][13] = -8'd21;
        rom[190][14] = -8'd16;
        rom[190][15] = 8'd29;
        rom[190][16] = -8'd10;
        rom[190][17] = 8'd0;
        rom[190][18] = 8'd35;
        rom[190][19] = 8'd13;
        rom[190][20] = -8'd17;
        rom[190][21] = 8'd33;
        rom[190][22] = -8'd70;
        rom[190][23] = -8'd20;
        rom[190][24] = -8'd19;
        rom[190][25] = 8'd11;
        rom[190][26] = -8'd7;
        rom[190][27] = -8'd48;
        rom[190][28] = -8'd1;
        rom[190][29] = -8'd51;
        rom[190][30] = 8'd11;
        rom[190][31] = 8'd11;
        rom[190][32] = -8'd10;
        rom[190][33] = -8'd25;
        rom[190][34] = 8'd21;
        rom[190][35] = 8'd1;
        rom[190][36] = 8'd32;
        rom[190][37] = -8'd11;
        rom[190][38] = 8'd35;
        rom[190][39] = 8'd14;
        rom[190][40] = 8'd21;
        rom[190][41] = 8'd27;
        rom[190][42] = -8'd46;
        rom[190][43] = -8'd45;
        rom[190][44] = -8'd2;
        rom[190][45] = 8'd3;
        rom[190][46] = -8'd28;
        rom[190][47] = -8'd4;
        rom[190][48] = -8'd58;
        rom[190][49] = -8'd8;
        rom[190][50] = 8'd7;
        rom[190][51] = 8'd23;
        rom[190][52] = 8'd2;
        rom[190][53] = -8'd19;
        rom[190][54] = -8'd19;
        rom[190][55] = -8'd12;
        rom[190][56] = 8'd12;
        rom[190][57] = -8'd30;
        rom[190][58] = -8'd10;
        rom[190][59] = -8'd56;
        rom[190][60] = -8'd8;
        rom[190][61] = -8'd36;
        rom[190][62] = 8'd2;
        rom[190][63] = -8'd15;
        rom[191][0] = -8'd30;
        rom[191][1] = -8'd5;
        rom[191][2] = -8'd24;
        rom[191][3] = 8'd2;
        rom[191][4] = -8'd24;
        rom[191][5] = -8'd11;
        rom[191][6] = -8'd9;
        rom[191][7] = 8'd14;
        rom[191][8] = -8'd31;
        rom[191][9] = -8'd34;
        rom[191][10] = 8'd54;
        rom[191][11] = 8'd19;
        rom[191][12] = -8'd15;
        rom[191][13] = -8'd14;
        rom[191][14] = -8'd47;
        rom[191][15] = -8'd4;
        rom[191][16] = 8'd3;
        rom[191][17] = -8'd9;
        rom[191][18] = 8'd15;
        rom[191][19] = -8'd1;
        rom[191][20] = -8'd1;
        rom[191][21] = 8'd9;
        rom[191][22] = 8'd0;
        rom[191][23] = -8'd8;
        rom[191][24] = 8'd9;
        rom[191][25] = -8'd80;
        rom[191][26] = -8'd11;
        rom[191][27] = -8'd40;
        rom[191][28] = -8'd57;
        rom[191][29] = -8'd56;
        rom[191][30] = 8'd11;
        rom[191][31] = -8'd20;
        rom[191][32] = -8'd49;
        rom[191][33] = -8'd3;
        rom[191][34] = 8'd19;
        rom[191][35] = -8'd13;
        rom[191][36] = -8'd2;
        rom[191][37] = 8'd19;
        rom[191][38] = 8'd48;
        rom[191][39] = -8'd21;
        rom[191][40] = 8'd10;
        rom[191][41] = 8'd33;
        rom[191][42] = -8'd18;
        rom[191][43] = 8'd6;
        rom[191][44] = -8'd40;
        rom[191][45] = 8'd13;
        rom[191][46] = 8'd14;
        rom[191][47] = 8'd5;
        rom[191][48] = -8'd22;
        rom[191][49] = 8'd9;
        rom[191][50] = -8'd1;
        rom[191][51] = -8'd21;
        rom[191][52] = -8'd6;
        rom[191][53] = -8'd12;
        rom[191][54] = 8'd24;
        rom[191][55] = -8'd12;
        rom[191][56] = 8'd8;
        rom[191][57] = 8'd17;
        rom[191][58] = 8'd6;
        rom[191][59] = 8'd46;
        rom[191][60] = -8'd98;
        rom[191][61] = 8'd56;
        rom[191][62] = -8'd53;
        rom[191][63] = -8'd18;
        rom[192][0] = -8'd13;
        rom[192][1] = 8'd1;
        rom[192][2] = -8'd28;
        rom[192][3] = -8'd17;
        rom[192][4] = -8'd35;
        rom[192][5] = 8'd11;
        rom[192][6] = 8'd7;
        rom[192][7] = -8'd6;
        rom[192][8] = -8'd34;
        rom[192][9] = 8'd34;
        rom[192][10] = 8'd1;
        rom[192][11] = 8'd8;
        rom[192][12] = -8'd8;
        rom[192][13] = -8'd11;
        rom[192][14] = 8'd10;
        rom[192][15] = 8'd6;
        rom[192][16] = 8'd21;
        rom[192][17] = -8'd44;
        rom[192][18] = -8'd1;
        rom[192][19] = -8'd9;
        rom[192][20] = -8'd8;
        rom[192][21] = -8'd34;
        rom[192][22] = 8'd14;
        rom[192][23] = -8'd25;
        rom[192][24] = 8'd17;
        rom[192][25] = -8'd12;
        rom[192][26] = -8'd24;
        rom[192][27] = -8'd20;
        rom[192][28] = -8'd23;
        rom[192][29] = 8'd8;
        rom[192][30] = -8'd7;
        rom[192][31] = -8'd27;
        rom[192][32] = -8'd12;
        rom[192][33] = -8'd18;
        rom[192][34] = -8'd31;
        rom[192][35] = -8'd30;
        rom[192][36] = -8'd34;
        rom[192][37] = 8'd25;
        rom[192][38] = -8'd15;
        rom[192][39] = -8'd12;
        rom[192][40] = -8'd28;
        rom[192][41] = -8'd81;
        rom[192][42] = 8'd16;
        rom[192][43] = 8'd3;
        rom[192][44] = -8'd21;
        rom[192][45] = 8'd31;
        rom[192][46] = 8'd3;
        rom[192][47] = 8'd30;
        rom[192][48] = -8'd33;
        rom[192][49] = -8'd3;
        rom[192][50] = -8'd2;
        rom[192][51] = -8'd58;
        rom[192][52] = 8'd11;
        rom[192][53] = -8'd31;
        rom[192][54] = 8'd2;
        rom[192][55] = 8'd22;
        rom[192][56] = -8'd25;
        rom[192][57] = 8'd3;
        rom[192][58] = -8'd1;
        rom[192][59] = 8'd34;
        rom[192][60] = 8'd15;
        rom[192][61] = -8'd50;
        rom[192][62] = 8'd14;
        rom[192][63] = 8'd7;
        rom[193][0] = -8'd37;
        rom[193][1] = -8'd44;
        rom[193][2] = -8'd9;
        rom[193][3] = -8'd5;
        rom[193][4] = -8'd8;
        rom[193][5] = -8'd18;
        rom[193][6] = -8'd100;
        rom[193][7] = -8'd41;
        rom[193][8] = 8'd13;
        rom[193][9] = -8'd11;
        rom[193][10] = -8'd88;
        rom[193][11] = -8'd68;
        rom[193][12] = 8'd30;
        rom[193][13] = -8'd20;
        rom[193][14] = 8'd0;
        rom[193][15] = -8'd39;
        rom[193][16] = -8'd41;
        rom[193][17] = 8'd34;
        rom[193][18] = -8'd31;
        rom[193][19] = 8'd4;
        rom[193][20] = -8'd8;
        rom[193][21] = -8'd2;
        rom[193][22] = 8'd13;
        rom[193][23] = -8'd67;
        rom[193][24] = 8'd19;
        rom[193][25] = -8'd40;
        rom[193][26] = 8'd1;
        rom[193][27] = 8'd7;
        rom[193][28] = 8'd6;
        rom[193][29] = -8'd55;
        rom[193][30] = 8'd0;
        rom[193][31] = -8'd32;
        rom[193][32] = -8'd2;
        rom[193][33] = -8'd56;
        rom[193][34] = -8'd2;
        rom[193][35] = 8'd24;
        rom[193][36] = -8'd7;
        rom[193][37] = -8'd23;
        rom[193][38] = -8'd27;
        rom[193][39] = 8'd21;
        rom[193][40] = 8'd26;
        rom[193][41] = -8'd13;
        rom[193][42] = 8'd4;
        rom[193][43] = -8'd13;
        rom[193][44] = -8'd12;
        rom[193][45] = -8'd2;
        rom[193][46] = -8'd50;
        rom[193][47] = 8'd45;
        rom[193][48] = 8'd28;
        rom[193][49] = 8'd20;
        rom[193][50] = -8'd3;
        rom[193][51] = 8'd16;
        rom[193][52] = -8'd13;
        rom[193][53] = -8'd40;
        rom[193][54] = 8'd37;
        rom[193][55] = -8'd44;
        rom[193][56] = 8'd48;
        rom[193][57] = 8'd16;
        rom[193][58] = -8'd63;
        rom[193][59] = 8'd4;
        rom[193][60] = -8'd32;
        rom[193][61] = -8'd5;
        rom[193][62] = -8'd28;
        rom[193][63] = -8'd20;
        rom[194][0] = 8'd3;
        rom[194][1] = -8'd9;
        rom[194][2] = -8'd47;
        rom[194][3] = 8'd9;
        rom[194][4] = -8'd41;
        rom[194][5] = -8'd30;
        rom[194][6] = -8'd64;
        rom[194][7] = 8'd13;
        rom[194][8] = -8'd25;
        rom[194][9] = 8'd23;
        rom[194][10] = 8'd53;
        rom[194][11] = 8'd0;
        rom[194][12] = 8'd29;
        rom[194][13] = 8'd13;
        rom[194][14] = -8'd48;
        rom[194][15] = 8'd9;
        rom[194][16] = -8'd47;
        rom[194][17] = 8'd7;
        rom[194][18] = 8'd10;
        rom[194][19] = 8'd4;
        rom[194][20] = -8'd5;
        rom[194][21] = -8'd13;
        rom[194][22] = 8'd8;
        rom[194][23] = 8'd13;
        rom[194][24] = -8'd27;
        rom[194][25] = -8'd1;
        rom[194][26] = 8'd12;
        rom[194][27] = -8'd10;
        rom[194][28] = 8'd5;
        rom[194][29] = 8'd3;
        rom[194][30] = 8'd12;
        rom[194][31] = -8'd45;
        rom[194][32] = -8'd44;
        rom[194][33] = -8'd48;
        rom[194][34] = -8'd9;
        rom[194][35] = 8'd0;
        rom[194][36] = -8'd45;
        rom[194][37] = -8'd3;
        rom[194][38] = 8'd13;
        rom[194][39] = -8'd13;
        rom[194][40] = -8'd33;
        rom[194][41] = 8'd7;
        rom[194][42] = -8'd19;
        rom[194][43] = -8'd57;
        rom[194][44] = -8'd28;
        rom[194][45] = -8'd5;
        rom[194][46] = 8'd65;
        rom[194][47] = -8'd28;
        rom[194][48] = 8'd26;
        rom[194][49] = -8'd23;
        rom[194][50] = -8'd8;
        rom[194][51] = 8'd19;
        rom[194][52] = -8'd17;
        rom[194][53] = -8'd54;
        rom[194][54] = 8'd7;
        rom[194][55] = -8'd18;
        rom[194][56] = -8'd26;
        rom[194][57] = -8'd18;
        rom[194][58] = -8'd11;
        rom[194][59] = 8'd3;
        rom[194][60] = -8'd76;
        rom[194][61] = -8'd9;
        rom[194][62] = -8'd8;
        rom[194][63] = -8'd37;
        rom[195][0] = -8'd32;
        rom[195][1] = 8'd24;
        rom[195][2] = -8'd4;
        rom[195][3] = -8'd8;
        rom[195][4] = 8'd26;
        rom[195][5] = -8'd9;
        rom[195][6] = 8'd31;
        rom[195][7] = 8'd25;
        rom[195][8] = -8'd1;
        rom[195][9] = -8'd21;
        rom[195][10] = 8'd12;
        rom[195][11] = -8'd19;
        rom[195][12] = -8'd7;
        rom[195][13] = -8'd1;
        rom[195][14] = -8'd5;
        rom[195][15] = 8'd27;
        rom[195][16] = -8'd41;
        rom[195][17] = -8'd39;
        rom[195][18] = 8'd22;
        rom[195][19] = 8'd22;
        rom[195][20] = -8'd11;
        rom[195][21] = -8'd35;
        rom[195][22] = -8'd1;
        rom[195][23] = 8'd9;
        rom[195][24] = -8'd2;
        rom[195][25] = 8'd9;
        rom[195][26] = -8'd7;
        rom[195][27] = 8'd22;
        rom[195][28] = -8'd3;
        rom[195][29] = 8'd27;
        rom[195][30] = -8'd27;
        rom[195][31] = -8'd13;
        rom[195][32] = -8'd3;
        rom[195][33] = -8'd25;
        rom[195][34] = -8'd12;
        rom[195][35] = -8'd9;
        rom[195][36] = 8'd48;
        rom[195][37] = 8'd39;
        rom[195][38] = -8'd12;
        rom[195][39] = 8'd32;
        rom[195][40] = -8'd27;
        rom[195][41] = 8'd4;
        rom[195][42] = 8'd19;
        rom[195][43] = 8'd5;
        rom[195][44] = 8'd5;
        rom[195][45] = -8'd25;
        rom[195][46] = 8'd30;
        rom[195][47] = -8'd47;
        rom[195][48] = 8'd22;
        rom[195][49] = 8'd6;
        rom[195][50] = -8'd33;
        rom[195][51] = -8'd33;
        rom[195][52] = 8'd27;
        rom[195][53] = -8'd10;
        rom[195][54] = -8'd16;
        rom[195][55] = -8'd14;
        rom[195][56] = 8'd1;
        rom[195][57] = -8'd84;
        rom[195][58] = -8'd17;
        rom[195][59] = -8'd8;
        rom[195][60] = 8'd8;
        rom[195][61] = 8'd1;
        rom[195][62] = 8'd23;
        rom[195][63] = 8'd40;
        rom[196][0] = -8'd8;
        rom[196][1] = -8'd21;
        rom[196][2] = 8'd20;
        rom[196][3] = -8'd8;
        rom[196][4] = -8'd5;
        rom[196][5] = -8'd13;
        rom[196][6] = -8'd24;
        rom[196][7] = -8'd10;
        rom[196][8] = -8'd1;
        rom[196][9] = -8'd5;
        rom[196][10] = -8'd16;
        rom[196][11] = -8'd18;
        rom[196][12] = -8'd58;
        rom[196][13] = -8'd8;
        rom[196][14] = 8'd6;
        rom[196][15] = 8'd26;
        rom[196][16] = -8'd9;
        rom[196][17] = 8'd16;
        rom[196][18] = 8'd30;
        rom[196][19] = -8'd6;
        rom[196][20] = -8'd9;
        rom[196][21] = -8'd45;
        rom[196][22] = -8'd13;
        rom[196][23] = 8'd37;
        rom[196][24] = -8'd22;
        rom[196][25] = -8'd13;
        rom[196][26] = -8'd12;
        rom[196][27] = 8'd16;
        rom[196][28] = -8'd15;
        rom[196][29] = 8'd6;
        rom[196][30] = 8'd0;
        rom[196][31] = -8'd13;
        rom[196][32] = 8'd19;
        rom[196][33] = 8'd20;
        rom[196][34] = -8'd43;
        rom[196][35] = -8'd16;
        rom[196][36] = -8'd48;
        rom[196][37] = -8'd15;
        rom[196][38] = -8'd41;
        rom[196][39] = 8'd24;
        rom[196][40] = -8'd25;
        rom[196][41] = -8'd44;
        rom[196][42] = 8'd14;
        rom[196][43] = 8'd6;
        rom[196][44] = 8'd4;
        rom[196][45] = -8'd22;
        rom[196][46] = -8'd54;
        rom[196][47] = -8'd26;
        rom[196][48] = 8'd0;
        rom[196][49] = -8'd10;
        rom[196][50] = -8'd11;
        rom[196][51] = -8'd15;
        rom[196][52] = 8'd2;
        rom[196][53] = -8'd27;
        rom[196][54] = 8'd28;
        rom[196][55] = -8'd7;
        rom[196][56] = 8'd1;
        rom[196][57] = -8'd10;
        rom[196][58] = 8'd30;
        rom[196][59] = 8'd11;
        rom[196][60] = -8'd8;
        rom[196][61] = 8'd5;
        rom[196][62] = 8'd7;
        rom[196][63] = -8'd7;
        rom[197][0] = 8'd6;
        rom[197][1] = -8'd11;
        rom[197][2] = 8'd1;
        rom[197][3] = -8'd1;
        rom[197][4] = -8'd6;
        rom[197][5] = 8'd1;
        rom[197][6] = -8'd9;
        rom[197][7] = -8'd5;
        rom[197][8] = 8'd0;
        rom[197][9] = -8'd7;
        rom[197][10] = 8'd5;
        rom[197][11] = -8'd1;
        rom[197][12] = 8'd8;
        rom[197][13] = -8'd4;
        rom[197][14] = 8'd4;
        rom[197][15] = 8'd4;
        rom[197][16] = 8'd0;
        rom[197][17] = -8'd5;
        rom[197][18] = -8'd10;
        rom[197][19] = 8'd8;
        rom[197][20] = -8'd1;
        rom[197][21] = -8'd2;
        rom[197][22] = 8'd9;
        rom[197][23] = 8'd10;
        rom[197][24] = 8'd17;
        rom[197][25] = 8'd11;
        rom[197][26] = 8'd3;
        rom[197][27] = -8'd1;
        rom[197][28] = -8'd11;
        rom[197][29] = -8'd5;
        rom[197][30] = 8'd11;
        rom[197][31] = -8'd1;
        rom[197][32] = -8'd13;
        rom[197][33] = 8'd10;
        rom[197][34] = 8'd0;
        rom[197][35] = 8'd9;
        rom[197][36] = 8'd2;
        rom[197][37] = 8'd12;
        rom[197][38] = 8'd12;
        rom[197][39] = 8'd5;
        rom[197][40] = 8'd4;
        rom[197][41] = 8'd0;
        rom[197][42] = 8'd4;
        rom[197][43] = -8'd1;
        rom[197][44] = 8'd0;
        rom[197][45] = -8'd1;
        rom[197][46] = -8'd1;
        rom[197][47] = 8'd7;
        rom[197][48] = -8'd5;
        rom[197][49] = -8'd3;
        rom[197][50] = -8'd3;
        rom[197][51] = -8'd8;
        rom[197][52] = 8'd5;
        rom[197][53] = 8'd12;
        rom[197][54] = -8'd4;
        rom[197][55] = 8'd7;
        rom[197][56] = -8'd6;
        rom[197][57] = 8'd9;
        rom[197][58] = 8'd1;
        rom[197][59] = 8'd4;
        rom[197][60] = 8'd1;
        rom[197][61] = 8'd8;
        rom[197][62] = 8'd1;
        rom[197][63] = -8'd11;
        rom[198][0] = -8'd11;
        rom[198][1] = -8'd59;
        rom[198][2] = -8'd12;
        rom[198][3] = 8'd6;
        rom[198][4] = -8'd6;
        rom[198][5] = 8'd20;
        rom[198][6] = -8'd35;
        rom[198][7] = -8'd6;
        rom[198][8] = 8'd0;
        rom[198][9] = 8'd43;
        rom[198][10] = -8'd7;
        rom[198][11] = 8'd6;
        rom[198][12] = 8'd16;
        rom[198][13] = -8'd19;
        rom[198][14] = -8'd13;
        rom[198][15] = -8'd38;
        rom[198][16] = -8'd24;
        rom[198][17] = -8'd19;
        rom[198][18] = -8'd41;
        rom[198][19] = 8'd9;
        rom[198][20] = -8'd11;
        rom[198][21] = -8'd95;
        rom[198][22] = 8'd11;
        rom[198][23] = -8'd12;
        rom[198][24] = 8'd5;
        rom[198][25] = 8'd0;
        rom[198][26] = 8'd15;
        rom[198][27] = 8'd36;
        rom[198][28] = 8'd4;
        rom[198][29] = 8'd1;
        rom[198][30] = -8'd72;
        rom[198][31] = -8'd15;
        rom[198][32] = -8'd32;
        rom[198][33] = 8'd10;
        rom[198][34] = 8'd12;
        rom[198][35] = 8'd20;
        rom[198][36] = 8'd7;
        rom[198][37] = -8'd22;
        rom[198][38] = 8'd8;
        rom[198][39] = -8'd33;
        rom[198][40] = 8'd18;
        rom[198][41] = -8'd20;
        rom[198][42] = 8'd4;
        rom[198][43] = -8'd2;
        rom[198][44] = 8'd22;
        rom[198][45] = -8'd20;
        rom[198][46] = -8'd20;
        rom[198][47] = -8'd84;
        rom[198][48] = -8'd49;
        rom[198][49] = 8'd3;
        rom[198][50] = 8'd17;
        rom[198][51] = 8'd3;
        rom[198][52] = -8'd15;
        rom[198][53] = 8'd23;
        rom[198][54] = -8'd10;
        rom[198][55] = 8'd52;
        rom[198][56] = -8'd3;
        rom[198][57] = 8'd35;
        rom[198][58] = -8'd5;
        rom[198][59] = -8'd3;
        rom[198][60] = -8'd14;
        rom[198][61] = -8'd27;
        rom[198][62] = -8'd39;
        rom[198][63] = 8'd7;
        rom[199][0] = -8'd22;
        rom[199][1] = 8'd8;
        rom[199][2] = -8'd29;
        rom[199][3] = -8'd16;
        rom[199][4] = -8'd46;
        rom[199][5] = 8'd6;
        rom[199][6] = -8'd3;
        rom[199][7] = -8'd25;
        rom[199][8] = 8'd4;
        rom[199][9] = 8'd0;
        rom[199][10] = 8'd7;
        rom[199][11] = -8'd23;
        rom[199][12] = -8'd22;
        rom[199][13] = 8'd13;
        rom[199][14] = -8'd25;
        rom[199][15] = -8'd23;
        rom[199][16] = -8'd7;
        rom[199][17] = 8'd1;
        rom[199][18] = -8'd5;
        rom[199][19] = 8'd21;
        rom[199][20] = -8'd5;
        rom[199][21] = 8'd18;
        rom[199][22] = -8'd33;
        rom[199][23] = 8'd18;
        rom[199][24] = 8'd31;
        rom[199][25] = 8'd3;
        rom[199][26] = -8'd30;
        rom[199][27] = 8'd6;
        rom[199][28] = 8'd21;
        rom[199][29] = -8'd16;
        rom[199][30] = -8'd1;
        rom[199][31] = -8'd16;
        rom[199][32] = 8'd9;
        rom[199][33] = 8'd32;
        rom[199][34] = 8'd14;
        rom[199][35] = 8'd27;
        rom[199][36] = -8'd8;
        rom[199][37] = -8'd32;
        rom[199][38] = 8'd13;
        rom[199][39] = 8'd6;
        rom[199][40] = 8'd8;
        rom[199][41] = 8'd21;
        rom[199][42] = 8'd6;
        rom[199][43] = 8'd3;
        rom[199][44] = 8'd23;
        rom[199][45] = 8'd74;
        rom[199][46] = 8'd23;
        rom[199][47] = 8'd18;
        rom[199][48] = -8'd13;
        rom[199][49] = 8'd8;
        rom[199][50] = -8'd9;
        rom[199][51] = -8'd11;
        rom[199][52] = 8'd20;
        rom[199][53] = -8'd16;
        rom[199][54] = 8'd44;
        rom[199][55] = -8'd17;
        rom[199][56] = 8'd32;
        rom[199][57] = 8'd8;
        rom[199][58] = -8'd50;
        rom[199][59] = 8'd8;
        rom[199][60] = -8'd17;
        rom[199][61] = -8'd33;
        rom[199][62] = -8'd22;
        rom[199][63] = 8'd50;
        rom[200][0] = -8'd30;
        rom[200][1] = 8'd6;
        rom[200][2] = -8'd22;
        rom[200][3] = -8'd11;
        rom[200][4] = 8'd15;
        rom[200][5] = -8'd27;
        rom[200][6] = -8'd22;
        rom[200][7] = -8'd30;
        rom[200][8] = 8'd7;
        rom[200][9] = -8'd2;
        rom[200][10] = 8'd13;
        rom[200][11] = -8'd63;
        rom[200][12] = 8'd24;
        rom[200][13] = -8'd20;
        rom[200][14] = 8'd8;
        rom[200][15] = 8'd7;
        rom[200][16] = -8'd3;
        rom[200][17] = -8'd40;
        rom[200][18] = 8'd24;
        rom[200][19] = -8'd8;
        rom[200][20] = -8'd5;
        rom[200][21] = 8'd5;
        rom[200][22] = -8'd31;
        rom[200][23] = -8'd20;
        rom[200][24] = -8'd7;
        rom[200][25] = 8'd15;
        rom[200][26] = -8'd17;
        rom[200][27] = -8'd18;
        rom[200][28] = -8'd1;
        rom[200][29] = -8'd5;
        rom[200][30] = -8'd40;
        rom[200][31] = -8'd24;
        rom[200][32] = 8'd16;
        rom[200][33] = 8'd5;
        rom[200][34] = -8'd13;
        rom[200][35] = -8'd39;
        rom[200][36] = 8'd19;
        rom[200][37] = -8'd10;
        rom[200][38] = -8'd29;
        rom[200][39] = 8'd4;
        rom[200][40] = -8'd35;
        rom[200][41] = -8'd31;
        rom[200][42] = -8'd23;
        rom[200][43] = 8'd23;
        rom[200][44] = 8'd31;
        rom[200][45] = -8'd14;
        rom[200][46] = -8'd10;
        rom[200][47] = -8'd6;
        rom[200][48] = -8'd36;
        rom[200][49] = 8'd8;
        rom[200][50] = 8'd1;
        rom[200][51] = -8'd15;
        rom[200][52] = 8'd24;
        rom[200][53] = 8'd24;
        rom[200][54] = 8'd12;
        rom[200][55] = 8'd25;
        rom[200][56] = -8'd30;
        rom[200][57] = 8'd10;
        rom[200][58] = -8'd12;
        rom[200][59] = -8'd28;
        rom[200][60] = -8'd11;
        rom[200][61] = -8'd24;
        rom[200][62] = -8'd11;
        rom[200][63] = -8'd19;
        rom[201][0] = -8'd10;
        rom[201][1] = 8'd10;
        rom[201][2] = 8'd15;
        rom[201][3] = -8'd68;
        rom[201][4] = 8'd42;
        rom[201][5] = 8'd5;
        rom[201][6] = -8'd10;
        rom[201][7] = 8'd20;
        rom[201][8] = -8'd31;
        rom[201][9] = 8'd31;
        rom[201][10] = 8'd12;
        rom[201][11] = -8'd13;
        rom[201][12] = -8'd33;
        rom[201][13] = 8'd5;
        rom[201][14] = 8'd21;
        rom[201][15] = -8'd32;
        rom[201][16] = 8'd7;
        rom[201][17] = 8'd1;
        rom[201][18] = 8'd9;
        rom[201][19] = -8'd71;
        rom[201][20] = -8'd16;
        rom[201][21] = -8'd32;
        rom[201][22] = -8'd34;
        rom[201][23] = 8'd10;
        rom[201][24] = 8'd3;
        rom[201][25] = -8'd6;
        rom[201][26] = 8'd19;
        rom[201][27] = -8'd63;
        rom[201][28] = -8'd4;
        rom[201][29] = -8'd26;
        rom[201][30] = -8'd48;
        rom[201][31] = 8'd40;
        rom[201][32] = -8'd23;
        rom[201][33] = 8'd5;
        rom[201][34] = 8'd23;
        rom[201][35] = -8'd40;
        rom[201][36] = 8'd2;
        rom[201][37] = 8'd38;
        rom[201][38] = 8'd13;
        rom[201][39] = -8'd16;
        rom[201][40] = -8'd9;
        rom[201][41] = -8'd30;
        rom[201][42] = -8'd58;
        rom[201][43] = -8'd23;
        rom[201][44] = 8'd35;
        rom[201][45] = -8'd27;
        rom[201][46] = -8'd10;
        rom[201][47] = -8'd5;
        rom[201][48] = -8'd36;
        rom[201][49] = -8'd24;
        rom[201][50] = -8'd58;
        rom[201][51] = 8'd14;
        rom[201][52] = 8'd21;
        rom[201][53] = 8'd10;
        rom[201][54] = -8'd47;
        rom[201][55] = 8'd16;
        rom[201][56] = -8'd8;
        rom[201][57] = -8'd3;
        rom[201][58] = -8'd9;
        rom[201][59] = 8'd26;
        rom[201][60] = 8'd16;
        rom[201][61] = 8'd18;
        rom[201][62] = 8'd34;
        rom[201][63] = 8'd0;
        rom[202][0] = 8'd19;
        rom[202][1] = -8'd46;
        rom[202][2] = 8'd1;
        rom[202][3] = 8'd12;
        rom[202][4] = -8'd14;
        rom[202][5] = -8'd4;
        rom[202][6] = 8'd37;
        rom[202][7] = -8'd8;
        rom[202][8] = -8'd2;
        rom[202][9] = -8'd6;
        rom[202][10] = -8'd1;
        rom[202][11] = 8'd16;
        rom[202][12] = -8'd4;
        rom[202][13] = 8'd31;
        rom[202][14] = -8'd46;
        rom[202][15] = 8'd21;
        rom[202][16] = -8'd36;
        rom[202][17] = -8'd36;
        rom[202][18] = -8'd45;
        rom[202][19] = -8'd1;
        rom[202][20] = -8'd2;
        rom[202][21] = -8'd1;
        rom[202][22] = -8'd5;
        rom[202][23] = -8'd39;
        rom[202][24] = 8'd0;
        rom[202][25] = -8'd15;
        rom[202][26] = 8'd5;
        rom[202][27] = 8'd15;
        rom[202][28] = -8'd67;
        rom[202][29] = -8'd14;
        rom[202][30] = 8'd17;
        rom[202][31] = 8'd24;
        rom[202][32] = 8'd42;
        rom[202][33] = -8'd13;
        rom[202][34] = -8'd42;
        rom[202][35] = 8'd4;
        rom[202][36] = -8'd14;
        rom[202][37] = 8'd37;
        rom[202][38] = 8'd43;
        rom[202][39] = -8'd18;
        rom[202][40] = 8'd4;
        rom[202][41] = -8'd10;
        rom[202][42] = 8'd13;
        rom[202][43] = -8'd15;
        rom[202][44] = 8'd8;
        rom[202][45] = 8'd25;
        rom[202][46] = -8'd7;
        rom[202][47] = -8'd2;
        rom[202][48] = -8'd23;
        rom[202][49] = 8'd24;
        rom[202][50] = -8'd17;
        rom[202][51] = 8'd27;
        rom[202][52] = 8'd7;
        rom[202][53] = -8'd42;
        rom[202][54] = -8'd37;
        rom[202][55] = 8'd11;
        rom[202][56] = 8'd2;
        rom[202][57] = -8'd11;
        rom[202][58] = 8'd17;
        rom[202][59] = 8'd12;
        rom[202][60] = 8'd30;
        rom[202][61] = -8'd13;
        rom[202][62] = -8'd41;
        rom[202][63] = 8'd6;
        rom[203][0] = 8'd1;
        rom[203][1] = 8'd14;
        rom[203][2] = 8'd20;
        rom[203][3] = -8'd14;
        rom[203][4] = -8'd2;
        rom[203][5] = 8'd2;
        rom[203][6] = 8'd3;
        rom[203][7] = -8'd7;
        rom[203][8] = 8'd46;
        rom[203][9] = 8'd19;
        rom[203][10] = -8'd22;
        rom[203][11] = 8'd7;
        rom[203][12] = -8'd10;
        rom[203][13] = 8'd43;
        rom[203][14] = -8'd37;
        rom[203][15] = -8'd6;
        rom[203][16] = 8'd2;
        rom[203][17] = -8'd11;
        rom[203][18] = -8'd3;
        rom[203][19] = -8'd16;
        rom[203][20] = -8'd6;
        rom[203][21] = -8'd6;
        rom[203][22] = 8'd4;
        rom[203][23] = 8'd30;
        rom[203][24] = -8'd17;
        rom[203][25] = 8'd5;
        rom[203][26] = 8'd19;
        rom[203][27] = -8'd19;
        rom[203][28] = 8'd16;
        rom[203][29] = 8'd1;
        rom[203][30] = -8'd10;
        rom[203][31] = -8'd17;
        rom[203][32] = -8'd63;
        rom[203][33] = 8'd22;
        rom[203][34] = 8'd17;
        rom[203][35] = 8'd18;
        rom[203][36] = -8'd25;
        rom[203][37] = 8'd16;
        rom[203][38] = -8'd25;
        rom[203][39] = -8'd18;
        rom[203][40] = -8'd8;
        rom[203][41] = 8'd27;
        rom[203][42] = -8'd69;
        rom[203][43] = 8'd13;
        rom[203][44] = -8'd20;
        rom[203][45] = -8'd2;
        rom[203][46] = -8'd26;
        rom[203][47] = 8'd10;
        rom[203][48] = -8'd40;
        rom[203][49] = -8'd8;
        rom[203][50] = -8'd19;
        rom[203][51] = -8'd4;
        rom[203][52] = -8'd33;
        rom[203][53] = -8'd11;
        rom[203][54] = 8'd17;
        rom[203][55] = -8'd20;
        rom[203][56] = 8'd5;
        rom[203][57] = -8'd24;
        rom[203][58] = -8'd29;
        rom[203][59] = 8'd19;
        rom[203][60] = -8'd28;
        rom[203][61] = -8'd8;
        rom[203][62] = -8'd5;
        rom[203][63] = 8'd15;
        rom[204][0] = 8'd0;
        rom[204][1] = 8'd50;
        rom[204][2] = 8'd51;
        rom[204][3] = 8'd35;
        rom[204][4] = 8'd6;
        rom[204][5] = -8'd1;
        rom[204][6] = 8'd0;
        rom[204][7] = -8'd69;
        rom[204][8] = 8'd14;
        rom[204][9] = -8'd7;
        rom[204][10] = 8'd8;
        rom[204][11] = 8'd15;
        rom[204][12] = -8'd12;
        rom[204][13] = 8'd12;
        rom[204][14] = 8'd23;
        rom[204][15] = -8'd5;
        rom[204][16] = -8'd1;
        rom[204][17] = -8'd31;
        rom[204][18] = 8'd16;
        rom[204][19] = -8'd5;
        rom[204][20] = 8'd0;
        rom[204][21] = -8'd21;
        rom[204][22] = 8'd16;
        rom[204][23] = -8'd30;
        rom[204][24] = -8'd55;
        rom[204][25] = 8'd32;
        rom[204][26] = -8'd1;
        rom[204][27] = -8'd33;
        rom[204][28] = -8'd11;
        rom[204][29] = 8'd8;
        rom[204][30] = 8'd32;
        rom[204][31] = -8'd13;
        rom[204][32] = 8'd24;
        rom[204][33] = 8'd23;
        rom[204][34] = 8'd20;
        rom[204][35] = -8'd9;
        rom[204][36] = 8'd25;
        rom[204][37] = -8'd33;
        rom[204][38] = 8'd6;
        rom[204][39] = 8'd35;
        rom[204][40] = -8'd59;
        rom[204][41] = -8'd13;
        rom[204][42] = -8'd49;
        rom[204][43] = 8'd11;
        rom[204][44] = 8'd24;
        rom[204][45] = -8'd4;
        rom[204][46] = 8'd45;
        rom[204][47] = 8'd46;
        rom[204][48] = 8'd12;
        rom[204][49] = -8'd5;
        rom[204][50] = 8'd42;
        rom[204][51] = 8'd15;
        rom[204][52] = -8'd23;
        rom[204][53] = -8'd21;
        rom[204][54] = 8'd69;
        rom[204][55] = 8'd25;
        rom[204][56] = -8'd7;
        rom[204][57] = -8'd29;
        rom[204][58] = -8'd33;
        rom[204][59] = -8'd4;
        rom[204][60] = 8'd6;
        rom[204][61] = -8'd19;
        rom[204][62] = 8'd13;
        rom[204][63] = 8'd33;
        rom[205][0] = -8'd2;
        rom[205][1] = 8'd2;
        rom[205][2] = -8'd43;
        rom[205][3] = -8'd8;
        rom[205][4] = 8'd27;
        rom[205][5] = 8'd36;
        rom[205][6] = 8'd42;
        rom[205][7] = 8'd20;
        rom[205][8] = 8'd14;
        rom[205][9] = 8'd16;
        rom[205][10] = 8'd2;
        rom[205][11] = 8'd1;
        rom[205][12] = -8'd11;
        rom[205][13] = 8'd5;
        rom[205][14] = -8'd61;
        rom[205][15] = -8'd4;
        rom[205][16] = 8'd28;
        rom[205][17] = -8'd25;
        rom[205][18] = 8'd0;
        rom[205][19] = 8'd11;
        rom[205][20] = -8'd1;
        rom[205][21] = 8'd12;
        rom[205][22] = -8'd22;
        rom[205][23] = 8'd12;
        rom[205][24] = -8'd4;
        rom[205][25] = -8'd13;
        rom[205][26] = 8'd24;
        rom[205][27] = -8'd4;
        rom[205][28] = -8'd6;
        rom[205][29] = 8'd20;
        rom[205][30] = -8'd27;
        rom[205][31] = -8'd14;
        rom[205][32] = -8'd6;
        rom[205][33] = 8'd8;
        rom[205][34] = -8'd59;
        rom[205][35] = -8'd33;
        rom[205][36] = -8'd4;
        rom[205][37] = 8'd7;
        rom[205][38] = -8'd26;
        rom[205][39] = 8'd17;
        rom[205][40] = -8'd12;
        rom[205][41] = -8'd8;
        rom[205][42] = 8'd0;
        rom[205][43] = -8'd16;
        rom[205][44] = 8'd4;
        rom[205][45] = 8'd21;
        rom[205][46] = -8'd18;
        rom[205][47] = -8'd7;
        rom[205][48] = -8'd17;
        rom[205][49] = -8'd30;
        rom[205][50] = -8'd19;
        rom[205][51] = -8'd32;
        rom[205][52] = 8'd3;
        rom[205][53] = -8'd5;
        rom[205][54] = 8'd5;
        rom[205][55] = 8'd2;
        rom[205][56] = -8'd21;
        rom[205][57] = -8'd9;
        rom[205][58] = 8'd1;
        rom[205][59] = -8'd38;
        rom[205][60] = 8'd5;
        rom[205][61] = -8'd1;
        rom[205][62] = -8'd32;
        rom[205][63] = -8'd1;
        rom[206][0] = -8'd23;
        rom[206][1] = -8'd2;
        rom[206][2] = 8'd21;
        rom[206][3] = 8'd0;
        rom[206][4] = 8'd17;
        rom[206][5] = -8'd11;
        rom[206][6] = 8'd2;
        rom[206][7] = -8'd49;
        rom[206][8] = 8'd18;
        rom[206][9] = -8'd30;
        rom[206][10] = 8'd3;
        rom[206][11] = 8'd26;
        rom[206][12] = -8'd24;
        rom[206][13] = -8'd11;
        rom[206][14] = -8'd13;
        rom[206][15] = -8'd23;
        rom[206][16] = -8'd59;
        rom[206][17] = -8'd33;
        rom[206][18] = 8'd24;
        rom[206][19] = 8'd20;
        rom[206][20] = -8'd8;
        rom[206][21] = 8'd40;
        rom[206][22] = -8'd20;
        rom[206][23] = 8'd24;
        rom[206][24] = -8'd44;
        rom[206][25] = 8'd53;
        rom[206][26] = 8'd4;
        rom[206][27] = 8'd8;
        rom[206][28] = -8'd10;
        rom[206][29] = 8'd23;
        rom[206][30] = 8'd14;
        rom[206][31] = 8'd4;
        rom[206][32] = 8'd19;
        rom[206][33] = 8'd29;
        rom[206][34] = 8'd20;
        rom[206][35] = -8'd20;
        rom[206][36] = 8'd42;
        rom[206][37] = -8'd8;
        rom[206][38] = -8'd33;
        rom[206][39] = -8'd27;
        rom[206][40] = -8'd12;
        rom[206][41] = -8'd4;
        rom[206][42] = -8'd35;
        rom[206][43] = -8'd4;
        rom[206][44] = -8'd22;
        rom[206][45] = -8'd13;
        rom[206][46] = -8'd11;
        rom[206][47] = -8'd79;
        rom[206][48] = -8'd27;
        rom[206][49] = -8'd22;
        rom[206][50] = -8'd2;
        rom[206][51] = -8'd5;
        rom[206][52] = 8'd41;
        rom[206][53] = 8'd21;
        rom[206][54] = -8'd12;
        rom[206][55] = -8'd32;
        rom[206][56] = -8'd3;
        rom[206][57] = 8'd8;
        rom[206][58] = 8'd16;
        rom[206][59] = -8'd12;
        rom[206][60] = -8'd23;
        rom[206][61] = 8'd17;
        rom[206][62] = 8'd36;
        rom[206][63] = -8'd10;
        rom[207][0] = -8'd5;
        rom[207][1] = -8'd57;
        rom[207][2] = -8'd24;
        rom[207][3] = 8'd15;
        rom[207][4] = -8'd52;
        rom[207][5] = 8'd9;
        rom[207][6] = -8'd26;
        rom[207][7] = -8'd19;
        rom[207][8] = -8'd23;
        rom[207][9] = -8'd23;
        rom[207][10] = -8'd25;
        rom[207][11] = 8'd0;
        rom[207][12] = -8'd12;
        rom[207][13] = 8'd5;
        rom[207][14] = -8'd3;
        rom[207][15] = -8'd30;
        rom[207][16] = 8'd5;
        rom[207][17] = 8'd57;
        rom[207][18] = 8'd24;
        rom[207][19] = 8'd3;
        rom[207][20] = -8'd18;
        rom[207][21] = -8'd2;
        rom[207][22] = -8'd22;
        rom[207][23] = 8'd17;
        rom[207][24] = 8'd1;
        rom[207][25] = -8'd22;
        rom[207][26] = 8'd9;
        rom[207][27] = -8'd16;
        rom[207][28] = -8'd24;
        rom[207][29] = 8'd9;
        rom[207][30] = -8'd11;
        rom[207][31] = -8'd10;
        rom[207][32] = 8'd26;
        rom[207][33] = 8'd6;
        rom[207][34] = 8'd21;
        rom[207][35] = 8'd38;
        rom[207][36] = 8'd26;
        rom[207][37] = 8'd23;
        rom[207][38] = 8'd12;
        rom[207][39] = 8'd8;
        rom[207][40] = -8'd31;
        rom[207][41] = -8'd9;
        rom[207][42] = -8'd11;
        rom[207][43] = -8'd17;
        rom[207][44] = -8'd16;
        rom[207][45] = -8'd12;
        rom[207][46] = 8'd14;
        rom[207][47] = -8'd16;
        rom[207][48] = 8'd15;
        rom[207][49] = -8'd11;
        rom[207][50] = -8'd10;
        rom[207][51] = 8'd18;
        rom[207][52] = 8'd1;
        rom[207][53] = -8'd22;
        rom[207][54] = 8'd18;
        rom[207][55] = -8'd121;
        rom[207][56] = -8'd9;
        rom[207][57] = -8'd30;
        rom[207][58] = 8'd21;
        rom[207][59] = -8'd1;
        rom[207][60] = 8'd0;
        rom[207][61] = 8'd19;
        rom[207][62] = -8'd9;
        rom[207][63] = -8'd21;
        rom[208][0] = 8'd10;
        rom[208][1] = -8'd9;
        rom[208][2] = 8'd2;
        rom[208][3] = -8'd7;
        rom[208][4] = 8'd4;
        rom[208][5] = 8'd3;
        rom[208][6] = 8'd4;
        rom[208][7] = -8'd9;
        rom[208][8] = -8'd7;
        rom[208][9] = 8'd4;
        rom[208][10] = 8'd8;
        rom[208][11] = 8'd2;
        rom[208][12] = -8'd6;
        rom[208][13] = -8'd4;
        rom[208][14] = -8'd4;
        rom[208][15] = -8'd6;
        rom[208][16] = 8'd6;
        rom[208][17] = 8'd1;
        rom[208][18] = -8'd8;
        rom[208][19] = 8'd7;
        rom[208][20] = -8'd6;
        rom[208][21] = 8'd8;
        rom[208][22] = -8'd1;
        rom[208][23] = 8'd2;
        rom[208][24] = -8'd7;
        rom[208][25] = 8'd5;
        rom[208][26] = 8'd9;
        rom[208][27] = -8'd4;
        rom[208][28] = 8'd3;
        rom[208][29] = -8'd7;
        rom[208][30] = -8'd3;
        rom[208][31] = -8'd7;
        rom[208][32] = 8'd7;
        rom[208][33] = 8'd1;
        rom[208][34] = -8'd6;
        rom[208][35] = -8'd1;
        rom[208][36] = -8'd1;
        rom[208][37] = 8'd8;
        rom[208][38] = 8'd0;
        rom[208][39] = -8'd4;
        rom[208][40] = -8'd6;
        rom[208][41] = 8'd2;
        rom[208][42] = -8'd6;
        rom[208][43] = 8'd8;
        rom[208][44] = 8'd2;
        rom[208][45] = 8'd3;
        rom[208][46] = -8'd7;
        rom[208][47] = 8'd1;
        rom[208][48] = -8'd2;
        rom[208][49] = 8'd4;
        rom[208][50] = 8'd4;
        rom[208][51] = 8'd8;
        rom[208][52] = 8'd4;
        rom[208][53] = 8'd8;
        rom[208][54] = 8'd6;
        rom[208][55] = 8'd2;
        rom[208][56] = 8'd3;
        rom[208][57] = -8'd4;
        rom[208][58] = 8'd10;
        rom[208][59] = 8'd9;
        rom[208][60] = -8'd5;
        rom[208][61] = -8'd7;
        rom[208][62] = -8'd1;
        rom[208][63] = -8'd8;
        rom[209][0] = -8'd9;
        rom[209][1] = 8'd5;
        rom[209][2] = -8'd79;
        rom[209][3] = -8'd30;
        rom[209][4] = -8'd1;
        rom[209][5] = 8'd12;
        rom[209][6] = 8'd36;
        rom[209][7] = -8'd11;
        rom[209][8] = 8'd20;
        rom[209][9] = 8'd38;
        rom[209][10] = 8'd11;
        rom[209][11] = -8'd11;
        rom[209][12] = -8'd29;
        rom[209][13] = 8'd23;
        rom[209][14] = 8'd31;
        rom[209][15] = 8'd54;
        rom[209][16] = 8'd6;
        rom[209][17] = -8'd36;
        rom[209][18] = -8'd15;
        rom[209][19] = -8'd16;
        rom[209][20] = -8'd4;
        rom[209][21] = -8'd33;
        rom[209][22] = -8'd37;
        rom[209][23] = -8'd36;
        rom[209][24] = 8'd26;
        rom[209][25] = -8'd29;
        rom[209][26] = -8'd14;
        rom[209][27] = 8'd68;
        rom[209][28] = -8'd47;
        rom[209][29] = 8'd30;
        rom[209][30] = -8'd17;
        rom[209][31] = 8'd6;
        rom[209][32] = 8'd5;
        rom[209][33] = 8'd11;
        rom[209][34] = -8'd25;
        rom[209][35] = -8'd25;
        rom[209][36] = -8'd52;
        rom[209][37] = 8'd33;
        rom[209][38] = -8'd8;
        rom[209][39] = 8'd8;
        rom[209][40] = 8'd0;
        rom[209][41] = 8'd11;
        rom[209][42] = -8'd1;
        rom[209][43] = 8'd17;
        rom[209][44] = 8'd8;
        rom[209][45] = 8'd8;
        rom[209][46] = -8'd5;
        rom[209][47] = -8'd15;
        rom[209][48] = -8'd37;
        rom[209][49] = 8'd6;
        rom[209][50] = 8'd6;
        rom[209][51] = 8'd6;
        rom[209][52] = 8'd20;
        rom[209][53] = 8'd20;
        rom[209][54] = 8'd13;
        rom[209][55] = 8'd5;
        rom[209][56] = -8'd12;
        rom[209][57] = 8'd2;
        rom[209][58] = 8'd17;
        rom[209][59] = -8'd40;
        rom[209][60] = 8'd16;
        rom[209][61] = -8'd18;
        rom[209][62] = -8'd26;
        rom[209][63] = -8'd7;
        rom[210][0] = -8'd34;
        rom[210][1] = 8'd23;
        rom[210][2] = -8'd29;
        rom[210][3] = -8'd38;
        rom[210][4] = -8'd21;
        rom[210][5] = -8'd6;
        rom[210][6] = 8'd17;
        rom[210][7] = -8'd13;
        rom[210][8] = 8'd21;
        rom[210][9] = 8'd5;
        rom[210][10] = 8'd33;
        rom[210][11] = -8'd28;
        rom[210][12] = -8'd17;
        rom[210][13] = -8'd32;
        rom[210][14] = 8'd26;
        rom[210][15] = 8'd7;
        rom[210][16] = -8'd33;
        rom[210][17] = -8'd16;
        rom[210][18] = -8'd57;
        rom[210][19] = -8'd2;
        rom[210][20] = -8'd3;
        rom[210][21] = 8'd7;
        rom[210][22] = -8'd7;
        rom[210][23] = -8'd28;
        rom[210][24] = -8'd2;
        rom[210][25] = -8'd16;
        rom[210][26] = -8'd68;
        rom[210][27] = 8'd10;
        rom[210][28] = 8'd26;
        rom[210][29] = 8'd9;
        rom[210][30] = -8'd35;
        rom[210][31] = 8'd12;
        rom[210][32] = 8'd7;
        rom[210][33] = 8'd13;
        rom[210][34] = -8'd13;
        rom[210][35] = -8'd15;
        rom[210][36] = -8'd16;
        rom[210][37] = -8'd1;
        rom[210][38] = -8'd66;
        rom[210][39] = 8'd20;
        rom[210][40] = -8'd5;
        rom[210][41] = 8'd3;
        rom[210][42] = -8'd28;
        rom[210][43] = -8'd40;
        rom[210][44] = 8'd6;
        rom[210][45] = -8'd6;
        rom[210][46] = 8'd11;
        rom[210][47] = -8'd58;
        rom[210][48] = -8'd29;
        rom[210][49] = -8'd27;
        rom[210][50] = -8'd17;
        rom[210][51] = -8'd14;
        rom[210][52] = -8'd36;
        rom[210][53] = -8'd29;
        rom[210][54] = -8'd5;
        rom[210][55] = 8'd50;
        rom[210][56] = 8'd3;
        rom[210][57] = -8'd33;
        rom[210][58] = -8'd34;
        rom[210][59] = -8'd43;
        rom[210][60] = -8'd18;
        rom[210][61] = 8'd18;
        rom[210][62] = 8'd19;
        rom[210][63] = 8'd24;
        rom[211][0] = -8'd67;
        rom[211][1] = -8'd43;
        rom[211][2] = -8'd2;
        rom[211][3] = -8'd42;
        rom[211][4] = 8'd1;
        rom[211][5] = -8'd13;
        rom[211][6] = -8'd43;
        rom[211][7] = -8'd20;
        rom[211][8] = -8'd33;
        rom[211][9] = 8'd11;
        rom[211][10] = -8'd27;
        rom[211][11] = -8'd45;
        rom[211][12] = -8'd22;
        rom[211][13] = -8'd2;
        rom[211][14] = -8'd4;
        rom[211][15] = 8'd0;
        rom[211][16] = -8'd10;
        rom[211][17] = -8'd17;
        rom[211][18] = -8'd47;
        rom[211][19] = -8'd78;
        rom[211][20] = 8'd0;
        rom[211][21] = -8'd26;
        rom[211][22] = -8'd26;
        rom[211][23] = -8'd71;
        rom[211][24] = -8'd29;
        rom[211][25] = 8'd15;
        rom[211][26] = -8'd24;
        rom[211][27] = -8'd61;
        rom[211][28] = -8'd11;
        rom[211][29] = 8'd12;
        rom[211][30] = -8'd19;
        rom[211][31] = 8'd25;
        rom[211][32] = -8'd55;
        rom[211][33] = 8'd9;
        rom[211][34] = -8'd4;
        rom[211][35] = 8'd9;
        rom[211][36] = -8'd39;
        rom[211][37] = -8'd8;
        rom[211][38] = -8'd38;
        rom[211][39] = -8'd29;
        rom[211][40] = 8'd4;
        rom[211][41] = -8'd11;
        rom[211][42] = -8'd11;
        rom[211][43] = -8'd57;
        rom[211][44] = 8'd19;
        rom[211][45] = 8'd15;
        rom[211][46] = 8'd17;
        rom[211][47] = 8'd13;
        rom[211][48] = -8'd35;
        rom[211][49] = 8'd13;
        rom[211][50] = 8'd14;
        rom[211][51] = 8'd9;
        rom[211][52] = 8'd14;
        rom[211][53] = 8'd17;
        rom[211][54] = -8'd42;
        rom[211][55] = -8'd24;
        rom[211][56] = -8'd7;
        rom[211][57] = 8'd2;
        rom[211][58] = 8'd12;
        rom[211][59] = 8'd6;
        rom[211][60] = 8'd30;
        rom[211][61] = 8'd22;
        rom[211][62] = 8'd17;
        rom[211][63] = -8'd1;
        rom[212][0] = 8'd34;
        rom[212][1] = -8'd39;
        rom[212][2] = -8'd28;
        rom[212][3] = 8'd11;
        rom[212][4] = -8'd32;
        rom[212][5] = -8'd11;
        rom[212][6] = -8'd7;
        rom[212][7] = -8'd27;
        rom[212][8] = -8'd22;
        rom[212][9] = 8'd5;
        rom[212][10] = -8'd7;
        rom[212][11] = 8'd19;
        rom[212][12] = 8'd2;
        rom[212][13] = -8'd49;
        rom[212][14] = -8'd17;
        rom[212][15] = 8'd3;
        rom[212][16] = -8'd35;
        rom[212][17] = 8'd5;
        rom[212][18] = -8'd63;
        rom[212][19] = -8'd16;
        rom[212][20] = 8'd1;
        rom[212][21] = 8'd37;
        rom[212][22] = -8'd14;
        rom[212][23] = -8'd7;
        rom[212][24] = 8'd17;
        rom[212][25] = -8'd7;
        rom[212][26] = 8'd3;
        rom[212][27] = 8'd0;
        rom[212][28] = -8'd3;
        rom[212][29] = 8'd5;
        rom[212][30] = -8'd15;
        rom[212][31] = -8'd6;
        rom[212][32] = -8'd30;
        rom[212][33] = -8'd21;
        rom[212][34] = -8'd44;
        rom[212][35] = -8'd15;
        rom[212][36] = -8'd47;
        rom[212][37] = 8'd12;
        rom[212][38] = -8'd12;
        rom[212][39] = 8'd19;
        rom[212][40] = -8'd22;
        rom[212][41] = -8'd4;
        rom[212][42] = -8'd10;
        rom[212][43] = 8'd6;
        rom[212][44] = 8'd12;
        rom[212][45] = -8'd28;
        rom[212][46] = -8'd16;
        rom[212][47] = -8'd4;
        rom[212][48] = -8'd17;
        rom[212][49] = 8'd7;
        rom[212][50] = -8'd13;
        rom[212][51] = 8'd12;
        rom[212][52] = -8'd9;
        rom[212][53] = 8'd9;
        rom[212][54] = 8'd11;
        rom[212][55] = 8'd14;
        rom[212][56] = 8'd19;
        rom[212][57] = -8'd9;
        rom[212][58] = -8'd14;
        rom[212][59] = 8'd8;
        rom[212][60] = -8'd21;
        rom[212][61] = -8'd18;
        rom[212][62] = -8'd26;
        rom[212][63] = -8'd33;
        rom[213][0] = -8'd4;
        rom[213][1] = -8'd1;
        rom[213][2] = -8'd6;
        rom[213][3] = -8'd4;
        rom[213][4] = -8'd1;
        rom[213][5] = -8'd9;
        rom[213][6] = -8'd9;
        rom[213][7] = -8'd1;
        rom[213][8] = -8'd7;
        rom[213][9] = -8'd10;
        rom[213][10] = -8'd9;
        rom[213][11] = 8'd5;
        rom[213][12] = 8'd9;
        rom[213][13] = 8'd6;
        rom[213][14] = -8'd6;
        rom[213][15] = 8'd6;
        rom[213][16] = -8'd7;
        rom[213][17] = -8'd9;
        rom[213][18] = 8'd5;
        rom[213][19] = -8'd6;
        rom[213][20] = -8'd9;
        rom[213][21] = 8'd9;
        rom[213][22] = -8'd1;
        rom[213][23] = 8'd7;
        rom[213][24] = 8'd6;
        rom[213][25] = -8'd4;
        rom[213][26] = 8'd8;
        rom[213][27] = -8'd6;
        rom[213][28] = -8'd1;
        rom[213][29] = -8'd1;
        rom[213][30] = -8'd1;
        rom[213][31] = 8'd4;
        rom[213][32] = 8'd4;
        rom[213][33] = -8'd3;
        rom[213][34] = 8'd0;
        rom[213][35] = -8'd9;
        rom[213][36] = 8'd3;
        rom[213][37] = 8'd6;
        rom[213][38] = 8'd0;
        rom[213][39] = -8'd7;
        rom[213][40] = -8'd1;
        rom[213][41] = 8'd0;
        rom[213][42] = 8'd3;
        rom[213][43] = -8'd4;
        rom[213][44] = 8'd5;
        rom[213][45] = 8'd11;
        rom[213][46] = 8'd6;
        rom[213][47] = 8'd11;
        rom[213][48] = -8'd4;
        rom[213][49] = 8'd2;
        rom[213][50] = 8'd9;
        rom[213][51] = -8'd3;
        rom[213][52] = -8'd9;
        rom[213][53] = -8'd6;
        rom[213][54] = -8'd10;
        rom[213][55] = 8'd1;
        rom[213][56] = -8'd3;
        rom[213][57] = -8'd3;
        rom[213][58] = 8'd1;
        rom[213][59] = 8'd5;
        rom[213][60] = -8'd2;
        rom[213][61] = 8'd7;
        rom[213][62] = -8'd12;
        rom[213][63] = -8'd4;
        rom[214][0] = -8'd29;
        rom[214][1] = -8'd9;
        rom[214][2] = -8'd11;
        rom[214][3] = 8'd7;
        rom[214][4] = -8'd8;
        rom[214][5] = -8'd21;
        rom[214][6] = -8'd13;
        rom[214][7] = 8'd33;
        rom[214][8] = -8'd8;
        rom[214][9] = -8'd18;
        rom[214][10] = 8'd20;
        rom[214][11] = -8'd28;
        rom[214][12] = -8'd1;
        rom[214][13] = 8'd4;
        rom[214][14] = 8'd33;
        rom[214][15] = 8'd15;
        rom[214][16] = 8'd14;
        rom[214][17] = -8'd8;
        rom[214][18] = -8'd44;
        rom[214][19] = 8'd27;
        rom[214][20] = -8'd11;
        rom[214][21] = 8'd7;
        rom[214][22] = 8'd32;
        rom[214][23] = -8'd25;
        rom[214][24] = -8'd20;
        rom[214][25] = -8'd11;
        rom[214][26] = 8'd2;
        rom[214][27] = 8'd13;
        rom[214][28] = -8'd31;
        rom[214][29] = -8'd11;
        rom[214][30] = -8'd32;
        rom[214][31] = 8'd2;
        rom[214][32] = -8'd1;
        rom[214][33] = -8'd1;
        rom[214][34] = -8'd8;
        rom[214][35] = 8'd18;
        rom[214][36] = -8'd17;
        rom[214][37] = 8'd32;
        rom[214][38] = 8'd19;
        rom[214][39] = -8'd40;
        rom[214][40] = 8'd30;
        rom[214][41] = -8'd4;
        rom[214][42] = -8'd25;
        rom[214][43] = 8'd5;
        rom[214][44] = -8'd25;
        rom[214][45] = 8'd6;
        rom[214][46] = -8'd1;
        rom[214][47] = -8'd52;
        rom[214][48] = -8'd9;
        rom[214][49] = -8'd8;
        rom[214][50] = -8'd44;
        rom[214][51] = -8'd2;
        rom[214][52] = -8'd7;
        rom[214][53] = 8'd12;
        rom[214][54] = -8'd38;
        rom[214][55] = 8'd11;
        rom[214][56] = -8'd19;
        rom[214][57] = 8'd45;
        rom[214][58] = 8'd23;
        rom[214][59] = 8'd29;
        rom[214][60] = -8'd12;
        rom[214][61] = 8'd14;
        rom[214][62] = 8'd11;
        rom[214][63] = -8'd10;
        rom[215][0] = 8'd8;
        rom[215][1] = -8'd16;
        rom[215][2] = -8'd1;
        rom[215][3] = -8'd18;
        rom[215][4] = 8'd17;
        rom[215][5] = 8'd11;
        rom[215][6] = 8'd18;
        rom[215][7] = -8'd15;
        rom[215][8] = -8'd2;
        rom[215][9] = 8'd22;
        rom[215][10] = 8'd6;
        rom[215][11] = -8'd13;
        rom[215][12] = 8'd42;
        rom[215][13] = 8'd10;
        rom[215][14] = -8'd25;
        rom[215][15] = -8'd8;
        rom[215][16] = -8'd2;
        rom[215][17] = -8'd5;
        rom[215][18] = 8'd31;
        rom[215][19] = 8'd4;
        rom[215][20] = 8'd0;
        rom[215][21] = -8'd9;
        rom[215][22] = -8'd12;
        rom[215][23] = -8'd1;
        rom[215][24] = 8'd6;
        rom[215][25] = 8'd18;
        rom[215][26] = -8'd4;
        rom[215][27] = -8'd23;
        rom[215][28] = 8'd18;
        rom[215][29] = 8'd3;
        rom[215][30] = -8'd16;
        rom[215][31] = 8'd18;
        rom[215][32] = -8'd2;
        rom[215][33] = -8'd50;
        rom[215][34] = -8'd5;
        rom[215][35] = -8'd5;
        rom[215][36] = -8'd27;
        rom[215][37] = -8'd12;
        rom[215][38] = -8'd11;
        rom[215][39] = -8'd7;
        rom[215][40] = 8'd14;
        rom[215][41] = -8'd5;
        rom[215][42] = -8'd14;
        rom[215][43] = 8'd13;
        rom[215][44] = -8'd29;
        rom[215][45] = 8'd19;
        rom[215][46] = -8'd8;
        rom[215][47] = 8'd65;
        rom[215][48] = -8'd2;
        rom[215][49] = -8'd17;
        rom[215][50] = -8'd9;
        rom[215][51] = -8'd27;
        rom[215][52] = 8'd23;
        rom[215][53] = 8'd6;
        rom[215][54] = -8'd7;
        rom[215][55] = 8'd17;
        rom[215][56] = 8'd31;
        rom[215][57] = -8'd11;
        rom[215][58] = -8'd6;
        rom[215][59] = -8'd36;
        rom[215][60] = -8'd3;
        rom[215][61] = 8'd10;
        rom[215][62] = -8'd26;
        rom[215][63] = -8'd1;
        rom[216][0] = 8'd29;
        rom[216][1] = 8'd8;
        rom[216][2] = -8'd1;
        rom[216][3] = 8'd2;
        rom[216][4] = -8'd10;
        rom[216][5] = 8'd25;
        rom[216][6] = -8'd18;
        rom[216][7] = 8'd17;
        rom[216][8] = 8'd15;
        rom[216][9] = -8'd7;
        rom[216][10] = 8'd23;
        rom[216][11] = -8'd23;
        rom[216][12] = 8'd17;
        rom[216][13] = 8'd13;
        rom[216][14] = -8'd24;
        rom[216][15] = 8'd14;
        rom[216][16] = 8'd5;
        rom[216][17] = -8'd36;
        rom[216][18] = 8'd19;
        rom[216][19] = 8'd39;
        rom[216][20] = 8'd3;
        rom[216][21] = -8'd15;
        rom[216][22] = -8'd1;
        rom[216][23] = 8'd33;
        rom[216][24] = -8'd45;
        rom[216][25] = -8'd40;
        rom[216][26] = 8'd34;
        rom[216][27] = 8'd6;
        rom[216][28] = 8'd33;
        rom[216][29] = -8'd5;
        rom[216][30] = -8'd11;
        rom[216][31] = 8'd4;
        rom[216][32] = 8'd25;
        rom[216][33] = 8'd30;
        rom[216][34] = -8'd12;
        rom[216][35] = 8'd49;
        rom[216][36] = -8'd20;
        rom[216][37] = 8'd9;
        rom[216][38] = -8'd3;
        rom[216][39] = -8'd3;
        rom[216][40] = -8'd17;
        rom[216][41] = 8'd30;
        rom[216][42] = 8'd19;
        rom[216][43] = -8'd9;
        rom[216][44] = -8'd18;
        rom[216][45] = 8'd7;
        rom[216][46] = 8'd35;
        rom[216][47] = -8'd19;
        rom[216][48] = 8'd26;
        rom[216][49] = 8'd10;
        rom[216][50] = 8'd14;
        rom[216][51] = -8'd41;
        rom[216][52] = 8'd30;
        rom[216][53] = 8'd3;
        rom[216][54] = 8'd11;
        rom[216][55] = -8'd18;
        rom[216][56] = 8'd8;
        rom[216][57] = 8'd5;
        rom[216][58] = -8'd31;
        rom[216][59] = -8'd14;
        rom[216][60] = -8'd4;
        rom[216][61] = 8'd24;
        rom[216][62] = -8'd48;
        rom[216][63] = -8'd9;
        rom[217][0] = 8'd1;
        rom[217][1] = -8'd18;
        rom[217][2] = -8'd12;
        rom[217][3] = 8'd2;
        rom[217][4] = -8'd29;
        rom[217][5] = 8'd3;
        rom[217][6] = 8'd2;
        rom[217][7] = 8'd1;
        rom[217][8] = 8'd7;
        rom[217][9] = 8'd14;
        rom[217][10] = 8'd18;
        rom[217][11] = -8'd26;
        rom[217][12] = 8'd40;
        rom[217][13] = -8'd32;
        rom[217][14] = 8'd2;
        rom[217][15] = -8'd4;
        rom[217][16] = -8'd20;
        rom[217][17] = 8'd12;
        rom[217][18] = -8'd7;
        rom[217][19] = 8'd3;
        rom[217][20] = -8'd2;
        rom[217][21] = -8'd3;
        rom[217][22] = 8'd7;
        rom[217][23] = -8'd1;
        rom[217][24] = 8'd22;
        rom[217][25] = 8'd35;
        rom[217][26] = 8'd32;
        rom[217][27] = 8'd34;
        rom[217][28] = -8'd48;
        rom[217][29] = -8'd2;
        rom[217][30] = 8'd41;
        rom[217][31] = 8'd7;
        rom[217][32] = 8'd7;
        rom[217][33] = -8'd18;
        rom[217][34] = -8'd10;
        rom[217][35] = -8'd39;
        rom[217][36] = 8'd50;
        rom[217][37] = -8'd11;
        rom[217][38] = -8'd19;
        rom[217][39] = -8'd3;
        rom[217][40] = -8'd25;
        rom[217][41] = 8'd10;
        rom[217][42] = 8'd15;
        rom[217][43] = 8'd13;
        rom[217][44] = 8'd31;
        rom[217][45] = -8'd7;
        rom[217][46] = 8'd22;
        rom[217][47] = -8'd43;
        rom[217][48] = -8'd42;
        rom[217][49] = -8'd34;
        rom[217][50] = 8'd10;
        rom[217][51] = 8'd37;
        rom[217][52] = -8'd20;
        rom[217][53] = 8'd7;
        rom[217][54] = -8'd12;
        rom[217][55] = -8'd49;
        rom[217][56] = -8'd12;
        rom[217][57] = -8'd21;
        rom[217][58] = -8'd6;
        rom[217][59] = -8'd4;
        rom[217][60] = -8'd11;
        rom[217][61] = -8'd56;
        rom[217][62] = 8'd1;
        rom[217][63] = 8'd2;
        rom[218][0] = -8'd2;
        rom[218][1] = -8'd25;
        rom[218][2] = 8'd41;
        rom[218][3] = 8'd14;
        rom[218][4] = 8'd18;
        rom[218][5] = 8'd55;
        rom[218][6] = 8'd52;
        rom[218][7] = -8'd11;
        rom[218][8] = 8'd3;
        rom[218][9] = 8'd24;
        rom[218][10] = 8'd15;
        rom[218][11] = -8'd3;
        rom[218][12] = -8'd72;
        rom[218][13] = -8'd7;
        rom[218][14] = -8'd21;
        rom[218][15] = -8'd21;
        rom[218][16] = 8'd11;
        rom[218][17] = 8'd13;
        rom[218][18] = 8'd2;
        rom[218][19] = -8'd3;
        rom[218][20] = 8'd3;
        rom[218][21] = -8'd19;
        rom[218][22] = -8'd20;
        rom[218][23] = -8'd37;
        rom[218][24] = -8'd6;
        rom[218][25] = 8'd10;
        rom[218][26] = -8'd3;
        rom[218][27] = -8'd9;
        rom[218][28] = -8'd21;
        rom[218][29] = -8'd76;
        rom[218][30] = -8'd62;
        rom[218][31] = -8'd31;
        rom[218][32] = 8'd17;
        rom[218][33] = 8'd28;
        rom[218][34] = 8'd13;
        rom[218][35] = -8'd11;
        rom[218][36] = 8'd16;
        rom[218][37] = -8'd4;
        rom[218][38] = 8'd24;
        rom[218][39] = -8'd15;
        rom[218][40] = 8'd6;
        rom[218][41] = 8'd9;
        rom[218][42] = 8'd9;
        rom[218][43] = -8'd50;
        rom[218][44] = 8'd22;
        rom[218][45] = 8'd20;
        rom[218][46] = -8'd10;
        rom[218][47] = -8'd8;
        rom[218][48] = 8'd23;
        rom[218][49] = -8'd54;
        rom[218][50] = 8'd13;
        rom[218][51] = 8'd22;
        rom[218][52] = 8'd4;
        rom[218][53] = 8'd1;
        rom[218][54] = -8'd7;
        rom[218][55] = 8'd13;
        rom[218][56] = 8'd24;
        rom[218][57] = 8'd9;
        rom[218][58] = -8'd68;
        rom[218][59] = 8'd28;
        rom[218][60] = 8'd17;
        rom[218][61] = 8'd20;
        rom[218][62] = -8'd17;
        rom[218][63] = -8'd19;
        rom[219][0] = 8'd34;
        rom[219][1] = -8'd15;
        rom[219][2] = 8'd13;
        rom[219][3] = -8'd13;
        rom[219][4] = -8'd10;
        rom[219][5] = -8'd4;
        rom[219][6] = -8'd51;
        rom[219][7] = -8'd10;
        rom[219][8] = 8'd20;
        rom[219][9] = 8'd15;
        rom[219][10] = -8'd45;
        rom[219][11] = -8'd25;
        rom[219][12] = 8'd6;
        rom[219][13] = -8'd8;
        rom[219][14] = 8'd22;
        rom[219][15] = -8'd7;
        rom[219][16] = 8'd19;
        rom[219][17] = 8'd33;
        rom[219][18] = 8'd42;
        rom[219][19] = -8'd2;
        rom[219][20] = -8'd6;
        rom[219][21] = 8'd3;
        rom[219][22] = 8'd11;
        rom[219][23] = 8'd7;
        rom[219][24] = 8'd6;
        rom[219][25] = -8'd1;
        rom[219][26] = 8'd12;
        rom[219][27] = 8'd33;
        rom[219][28] = -8'd9;
        rom[219][29] = 8'd7;
        rom[219][30] = 8'd15;
        rom[219][31] = 8'd10;
        rom[219][32] = -8'd1;
        rom[219][33] = 8'd49;
        rom[219][34] = -8'd49;
        rom[219][35] = 8'd3;
        rom[219][36] = 8'd5;
        rom[219][37] = 8'd42;
        rom[219][38] = 8'd11;
        rom[219][39] = 8'd6;
        rom[219][40] = -8'd3;
        rom[219][41] = 8'd11;
        rom[219][42] = 8'd29;
        rom[219][43] = -8'd26;
        rom[219][44] = -8'd3;
        rom[219][45] = 8'd39;
        rom[219][46] = 8'd54;
        rom[219][47] = 8'd34;
        rom[219][48] = 8'd45;
        rom[219][49] = -8'd9;
        rom[219][50] = 8'd6;
        rom[219][51] = -8'd4;
        rom[219][52] = 8'd9;
        rom[219][53] = 8'd8;
        rom[219][54] = -8'd3;
        rom[219][55] = 8'd25;
        rom[219][56] = 8'd4;
        rom[219][57] = -8'd2;
        rom[219][58] = 8'd1;
        rom[219][59] = 8'd46;
        rom[219][60] = -8'd9;
        rom[219][61] = -8'd14;
        rom[219][62] = -8'd1;
        rom[219][63] = 8'd8;
        rom[220][0] = -8'd64;
        rom[220][1] = -8'd11;
        rom[220][2] = -8'd30;
        rom[220][3] = -8'd6;
        rom[220][4] = 8'd11;
        rom[220][5] = -8'd21;
        rom[220][6] = -8'd11;
        rom[220][7] = 8'd15;
        rom[220][8] = -8'd1;
        rom[220][9] = 8'd18;
        rom[220][10] = 8'd16;
        rom[220][11] = 8'd30;
        rom[220][12] = -8'd71;
        rom[220][13] = -8'd14;
        rom[220][14] = -8'd11;
        rom[220][15] = -8'd8;
        rom[220][16] = -8'd14;
        rom[220][17] = -8'd7;
        rom[220][18] = 8'd13;
        rom[220][19] = -8'd52;
        rom[220][20] = -8'd4;
        rom[220][21] = -8'd52;
        rom[220][22] = -8'd42;
        rom[220][23] = -8'd25;
        rom[220][24] = -8'd30;
        rom[220][25] = 8'd16;
        rom[220][26] = 8'd6;
        rom[220][27] = 8'd40;
        rom[220][28] = 8'd19;
        rom[220][29] = -8'd41;
        rom[220][30] = 8'd19;
        rom[220][31] = 8'd28;
        rom[220][32] = -8'd59;
        rom[220][33] = -8'd58;
        rom[220][34] = 8'd34;
        rom[220][35] = -8'd4;
        rom[220][36] = -8'd19;
        rom[220][37] = -8'd1;
        rom[220][38] = -8'd42;
        rom[220][39] = -8'd30;
        rom[220][40] = 8'd2;
        rom[220][41] = -8'd23;
        rom[220][42] = -8'd30;
        rom[220][43] = 8'd24;
        rom[220][44] = 8'd32;
        rom[220][45] = 8'd22;
        rom[220][46] = 8'd1;
        rom[220][47] = -8'd14;
        rom[220][48] = -8'd13;
        rom[220][49] = 8'd29;
        rom[220][50] = 8'd3;
        rom[220][51] = 8'd39;
        rom[220][52] = 8'd18;
        rom[220][53] = 8'd9;
        rom[220][54] = -8'd2;
        rom[220][55] = -8'd35;
        rom[220][56] = 8'd20;
        rom[220][57] = 8'd13;
        rom[220][58] = 8'd3;
        rom[220][59] = -8'd26;
        rom[220][60] = 8'd3;
        rom[220][61] = 8'd22;
        rom[220][62] = -8'd15;
        rom[220][63] = -8'd8;
        rom[221][0] = 8'd53;
        rom[221][1] = -8'd71;
        rom[221][2] = 8'd13;
        rom[221][3] = 8'd12;
        rom[221][4] = -8'd9;
        rom[221][5] = -8'd13;
        rom[221][6] = -8'd33;
        rom[221][7] = -8'd9;
        rom[221][8] = -8'd26;
        rom[221][9] = 8'd17;
        rom[221][10] = 8'd49;
        rom[221][11] = 8'd8;
        rom[221][12] = -8'd40;
        rom[221][13] = 8'd54;
        rom[221][14] = -8'd10;
        rom[221][15] = -8'd20;
        rom[221][16] = 8'd31;
        rom[221][17] = 8'd2;
        rom[221][18] = -8'd2;
        rom[221][19] = -8'd6;
        rom[221][20] = -8'd4;
        rom[221][21] = 8'd12;
        rom[221][22] = 8'd26;
        rom[221][23] = -8'd27;
        rom[221][24] = -8'd48;
        rom[221][25] = 8'd19;
        rom[221][26] = 8'd17;
        rom[221][27] = -8'd71;
        rom[221][28] = -8'd28;
        rom[221][29] = -8'd24;
        rom[221][30] = -8'd7;
        rom[221][31] = 8'd30;
        rom[221][32] = -8'd20;
        rom[221][33] = 8'd13;
        rom[221][34] = 8'd6;
        rom[221][35] = 8'd12;
        rom[221][36] = -8'd9;
        rom[221][37] = -8'd10;
        rom[221][38] = -8'd30;
        rom[221][39] = -8'd54;
        rom[221][40] = -8'd6;
        rom[221][41] = -8'd2;
        rom[221][42] = -8'd38;
        rom[221][43] = -8'd23;
        rom[221][44] = 8'd11;
        rom[221][45] = 8'd15;
        rom[221][46] = 8'd18;
        rom[221][47] = 8'd16;
        rom[221][48] = -8'd32;
        rom[221][49] = -8'd20;
        rom[221][50] = 8'd22;
        rom[221][51] = 8'd9;
        rom[221][52] = 8'd5;
        rom[221][53] = -8'd10;
        rom[221][54] = -8'd56;
        rom[221][55] = -8'd13;
        rom[221][56] = 8'd5;
        rom[221][57] = 8'd11;
        rom[221][58] = 8'd5;
        rom[221][59] = -8'd58;
        rom[221][60] = -8'd71;
        rom[221][61] = -8'd37;
        rom[221][62] = 8'd7;
        rom[221][63] = 8'd17;
        rom[222][0] = 8'd1;
        rom[222][1] = 8'd0;
        rom[222][2] = -8'd33;
        rom[222][3] = -8'd29;
        rom[222][4] = 8'd26;
        rom[222][5] = -8'd13;
        rom[222][6] = -8'd5;
        rom[222][7] = -8'd46;
        rom[222][8] = 8'd23;
        rom[222][9] = 8'd23;
        rom[222][10] = -8'd9;
        rom[222][11] = 8'd2;
        rom[222][12] = -8'd1;
        rom[222][13] = -8'd14;
        rom[222][14] = -8'd48;
        rom[222][15] = -8'd15;
        rom[222][16] = 8'd32;
        rom[222][17] = 8'd11;
        rom[222][18] = -8'd46;
        rom[222][19] = -8'd20;
        rom[222][20] = 8'd0;
        rom[222][21] = 8'd21;
        rom[222][22] = 8'd5;
        rom[222][23] = -8'd11;
        rom[222][24] = 8'd7;
        rom[222][25] = -8'd107;
        rom[222][26] = 8'd11;
        rom[222][27] = -8'd26;
        rom[222][28] = -8'd33;
        rom[222][29] = -8'd26;
        rom[222][30] = -8'd1;
        rom[222][31] = -8'd11;
        rom[222][32] = -8'd15;
        rom[222][33] = -8'd28;
        rom[222][34] = -8'd47;
        rom[222][35] = 8'd8;
        rom[222][36] = -8'd20;
        rom[222][37] = 8'd17;
        rom[222][38] = 8'd6;
        rom[222][39] = 8'd35;
        rom[222][40] = -8'd11;
        rom[222][41] = 8'd13;
        rom[222][42] = -8'd37;
        rom[222][43] = -8'd16;
        rom[222][44] = -8'd46;
        rom[222][45] = -8'd18;
        rom[222][46] = -8'd21;
        rom[222][47] = 8'd20;
        rom[222][48] = -8'd7;
        rom[222][49] = -8'd12;
        rom[222][50] = -8'd18;
        rom[222][51] = -8'd34;
        rom[222][52] = -8'd15;
        rom[222][53] = -8'd54;
        rom[222][54] = -8'd15;
        rom[222][55] = 8'd30;
        rom[222][56] = 8'd19;
        rom[222][57] = 8'd2;
        rom[222][58] = -8'd12;
        rom[222][59] = 8'd2;
        rom[222][60] = 8'd22;
        rom[222][61] = 8'd2;
        rom[222][62] = -8'd5;
        rom[222][63] = 8'd6;
        rom[223][0] = 8'd18;
        rom[223][1] = -8'd50;
        rom[223][2] = -8'd2;
        rom[223][3] = -8'd16;
        rom[223][4] = -8'd5;
        rom[223][5] = -8'd55;
        rom[223][6] = 8'd2;
        rom[223][7] = -8'd9;
        rom[223][8] = -8'd18;
        rom[223][9] = 8'd4;
        rom[223][10] = 8'd15;
        rom[223][11] = -8'd63;
        rom[223][12] = 8'd12;
        rom[223][13] = -8'd54;
        rom[223][14] = 8'd11;
        rom[223][15] = 8'd5;
        rom[223][16] = -8'd12;
        rom[223][17] = 8'd8;
        rom[223][18] = -8'd30;
        rom[223][19] = -8'd26;
        rom[223][20] = -8'd16;
        rom[223][21] = -8'd72;
        rom[223][22] = -8'd21;
        rom[223][23] = -8'd56;
        rom[223][24] = 8'd5;
        rom[223][25] = 8'd12;
        rom[223][26] = -8'd4;
        rom[223][27] = -8'd12;
        rom[223][28] = -8'd12;
        rom[223][29] = 8'd5;
        rom[223][30] = -8'd26;
        rom[223][31] = -8'd1;
        rom[223][32] = -8'd34;
        rom[223][33] = 8'd35;
        rom[223][34] = -8'd2;
        rom[223][35] = -8'd31;
        rom[223][36] = -8'd6;
        rom[223][37] = 8'd8;
        rom[223][38] = -8'd9;
        rom[223][39] = 8'd1;
        rom[223][40] = -8'd47;
        rom[223][41] = 8'd16;
        rom[223][42] = 8'd20;
        rom[223][43] = -8'd49;
        rom[223][44] = 8'd1;
        rom[223][45] = -8'd40;
        rom[223][46] = -8'd11;
        rom[223][47] = -8'd10;
        rom[223][48] = -8'd20;
        rom[223][49] = -8'd54;
        rom[223][50] = 8'd9;
        rom[223][51] = -8'd10;
        rom[223][52] = -8'd9;
        rom[223][53] = -8'd4;
        rom[223][54] = -8'd11;
        rom[223][55] = -8'd18;
        rom[223][56] = -8'd21;
        rom[223][57] = 8'd14;
        rom[223][58] = 8'd2;
        rom[223][59] = 8'd7;
        rom[223][60] = 8'd18;
        rom[223][61] = 8'd7;
        rom[223][62] = -8'd14;
        rom[223][63] = 8'd26;
        rom[224][0] = -8'd5;
        rom[224][1] = 8'd32;
        rom[224][2] = 8'd5;
        rom[224][3] = 8'd13;
        rom[224][4] = 8'd1;
        rom[224][5] = 8'd3;
        rom[224][6] = -8'd8;
        rom[224][7] = 8'd16;
        rom[224][8] = 8'd0;
        rom[224][9] = -8'd38;
        rom[224][10] = -8'd37;
        rom[224][11] = -8'd19;
        rom[224][12] = -8'd13;
        rom[224][13] = -8'd46;
        rom[224][14] = 8'd0;
        rom[224][15] = -8'd32;
        rom[224][16] = -8'd51;
        rom[224][17] = -8'd10;
        rom[224][18] = -8'd9;
        rom[224][19] = 8'd3;
        rom[224][20] = -8'd13;
        rom[224][21] = -8'd11;
        rom[224][22] = -8'd1;
        rom[224][23] = 8'd18;
        rom[224][24] = -8'd14;
        rom[224][25] = -8'd25;
        rom[224][26] = -8'd22;
        rom[224][27] = 8'd37;
        rom[224][28] = -8'd27;
        rom[224][29] = 8'd11;
        rom[224][30] = -8'd46;
        rom[224][31] = -8'd25;
        rom[224][32] = 8'd4;
        rom[224][33] = -8'd25;
        rom[224][34] = -8'd23;
        rom[224][35] = 8'd10;
        rom[224][36] = -8'd26;
        rom[224][37] = -8'd9;
        rom[224][38] = -8'd38;
        rom[224][39] = -8'd26;
        rom[224][40] = 8'd17;
        rom[224][41] = -8'd11;
        rom[224][42] = -8'd12;
        rom[224][43] = -8'd15;
        rom[224][44] = -8'd9;
        rom[224][45] = -8'd3;
        rom[224][46] = 8'd15;
        rom[224][47] = -8'd57;
        rom[224][48] = 8'd36;
        rom[224][49] = 8'd18;
        rom[224][50] = 8'd14;
        rom[224][51] = 8'd14;
        rom[224][52] = -8'd1;
        rom[224][53] = -8'd14;
        rom[224][54] = 8'd25;
        rom[224][55] = -8'd33;
        rom[224][56] = -8'd9;
        rom[224][57] = -8'd16;
        rom[224][58] = 8'd5;
        rom[224][59] = 8'd21;
        rom[224][60] = -8'd5;
        rom[224][61] = 8'd10;
        rom[224][62] = 8'd21;
        rom[224][63] = -8'd19;
        rom[225][0] = 8'd42;
        rom[225][1] = -8'd31;
        rom[225][2] = -8'd7;
        rom[225][3] = 8'd25;
        rom[225][4] = 8'd12;
        rom[225][5] = -8'd16;
        rom[225][6] = 8'd9;
        rom[225][7] = 8'd11;
        rom[225][8] = 8'd0;
        rom[225][9] = -8'd25;
        rom[225][10] = 8'd34;
        rom[225][11] = 8'd24;
        rom[225][12] = 8'd1;
        rom[225][13] = -8'd28;
        rom[225][14] = -8'd80;
        rom[225][15] = 8'd41;
        rom[225][16] = 8'd21;
        rom[225][17] = 8'd14;
        rom[225][18] = 8'd3;
        rom[225][19] = -8'd21;
        rom[225][20] = -8'd5;
        rom[225][21] = -8'd14;
        rom[225][22] = -8'd12;
        rom[225][23] = 8'd9;
        rom[225][24] = -8'd13;
        rom[225][25] = 8'd33;
        rom[225][26] = 8'd14;
        rom[225][27] = -8'd26;
        rom[225][28] = 8'd16;
        rom[225][29] = -8'd4;
        rom[225][30] = -8'd7;
        rom[225][31] = 8'd4;
        rom[225][32] = 8'd30;
        rom[225][33] = 8'd32;
        rom[225][34] = -8'd55;
        rom[225][35] = 8'd4;
        rom[225][36] = 8'd5;
        rom[225][37] = 8'd12;
        rom[225][38] = -8'd14;
        rom[225][39] = 8'd8;
        rom[225][40] = -8'd18;
        rom[225][41] = -8'd26;
        rom[225][42] = 8'd12;
        rom[225][43] = -8'd30;
        rom[225][44] = 8'd11;
        rom[225][45] = 8'd35;
        rom[225][46] = 8'd40;
        rom[225][47] = -8'd43;
        rom[225][48] = -8'd49;
        rom[225][49] = -8'd8;
        rom[225][50] = 8'd28;
        rom[225][51] = 8'd17;
        rom[225][52] = -8'd68;
        rom[225][53] = -8'd7;
        rom[225][54] = 8'd25;
        rom[225][55] = -8'd7;
        rom[225][56] = -8'd37;
        rom[225][57] = 8'd2;
        rom[225][58] = -8'd29;
        rom[225][59] = 8'd23;
        rom[225][60] = -8'd3;
        rom[225][61] = 8'd2;
        rom[225][62] = 8'd39;
        rom[225][63] = -8'd37;
        rom[226][0] = -8'd11;
        rom[226][1] = 8'd27;
        rom[226][2] = 8'd35;
        rom[226][3] = -8'd17;
        rom[226][4] = -8'd6;
        rom[226][5] = 8'd10;
        rom[226][6] = 8'd17;
        rom[226][7] = 8'd20;
        rom[226][8] = 8'd14;
        rom[226][9] = 8'd24;
        rom[226][10] = 8'd7;
        rom[226][11] = 8'd22;
        rom[226][12] = -8'd37;
        rom[226][13] = -8'd18;
        rom[226][14] = 8'd26;
        rom[226][15] = -8'd2;
        rom[226][16] = -8'd2;
        rom[226][17] = -8'd7;
        rom[226][18] = 8'd1;
        rom[226][19] = -8'd32;
        rom[226][20] = -8'd1;
        rom[226][21] = -8'd2;
        rom[226][22] = 8'd14;
        rom[226][23] = 8'd36;
        rom[226][24] = 8'd18;
        rom[226][25] = -8'd8;
        rom[226][26] = 8'd33;
        rom[226][27] = -8'd90;
        rom[226][28] = -8'd14;
        rom[226][29] = -8'd27;
        rom[226][30] = -8'd8;
        rom[226][31] = -8'd20;
        rom[226][32] = 8'd6;
        rom[226][33] = -8'd29;
        rom[226][34] = 8'd3;
        rom[226][35] = 8'd1;
        rom[226][36] = 8'd26;
        rom[226][37] = -8'd8;
        rom[226][38] = 8'd9;
        rom[226][39] = 8'd29;
        rom[226][40] = 8'd16;
        rom[226][41] = -8'd29;
        rom[226][42] = -8'd24;
        rom[226][43] = -8'd43;
        rom[226][44] = -8'd7;
        rom[226][45] = -8'd5;
        rom[226][46] = -8'd15;
        rom[226][47] = -8'd28;
        rom[226][48] = 8'd21;
        rom[226][49] = 8'd40;
        rom[226][50] = 8'd13;
        rom[226][51] = 8'd23;
        rom[226][52] = 8'd13;
        rom[226][53] = 8'd3;
        rom[226][54] = -8'd13;
        rom[226][55] = 8'd0;
        rom[226][56] = -8'd23;
        rom[226][57] = -8'd12;
        rom[226][58] = -8'd57;
        rom[226][59] = 8'd26;
        rom[226][60] = -8'd7;
        rom[226][61] = 8'd43;
        rom[226][62] = -8'd11;
        rom[226][63] = 8'd14;
        rom[227][0] = -8'd9;
        rom[227][1] = -8'd3;
        rom[227][2] = -8'd5;
        rom[227][3] = -8'd55;
        rom[227][4] = -8'd33;
        rom[227][5] = -8'd12;
        rom[227][6] = -8'd4;
        rom[227][7] = -8'd18;
        rom[227][8] = 8'd19;
        rom[227][9] = 8'd7;
        rom[227][10] = -8'd30;
        rom[227][11] = 8'd17;
        rom[227][12] = -8'd47;
        rom[227][13] = -8'd15;
        rom[227][14] = -8'd3;
        rom[227][15] = -8'd18;
        rom[227][16] = 8'd50;
        rom[227][17] = -8'd15;
        rom[227][18] = -8'd42;
        rom[227][19] = -8'd49;
        rom[227][20] = 8'd2;
        rom[227][21] = -8'd48;
        rom[227][22] = -8'd10;
        rom[227][23] = -8'd8;
        rom[227][24] = -8'd14;
        rom[227][25] = 8'd19;
        rom[227][26] = -8'd62;
        rom[227][27] = -8'd6;
        rom[227][28] = 8'd0;
        rom[227][29] = 8'd15;
        rom[227][30] = -8'd37;
        rom[227][31] = 8'd1;
        rom[227][32] = -8'd32;
        rom[227][33] = -8'd6;
        rom[227][34] = -8'd7;
        rom[227][35] = 8'd12;
        rom[227][36] = -8'd3;
        rom[227][37] = -8'd1;
        rom[227][38] = -8'd35;
        rom[227][39] = -8'd19;
        rom[227][40] = -8'd18;
        rom[227][41] = -8'd21;
        rom[227][42] = -8'd79;
        rom[227][43] = 8'd6;
        rom[227][44] = 8'd3;
        rom[227][45] = -8'd20;
        rom[227][46] = -8'd45;
        rom[227][47] = 8'd8;
        rom[227][48] = -8'd60;
        rom[227][49] = 8'd22;
        rom[227][50] = -8'd6;
        rom[227][51] = 8'd15;
        rom[227][52] = -8'd39;
        rom[227][53] = -8'd11;
        rom[227][54] = 8'd7;
        rom[227][55] = -8'd15;
        rom[227][56] = -8'd14;
        rom[227][57] = -8'd5;
        rom[227][58] = 8'd18;
        rom[227][59] = 8'd15;
        rom[227][60] = -8'd36;
        rom[227][61] = -8'd25;
        rom[227][62] = -8'd12;
        rom[227][63] = 8'd24;
        rom[228][0] = -8'd4;
        rom[228][1] = -8'd7;
        rom[228][2] = -8'd5;
        rom[228][3] = -8'd19;
        rom[228][4] = -8'd7;
        rom[228][5] = -8'd23;
        rom[228][6] = 8'd8;
        rom[228][7] = -8'd40;
        rom[228][8] = -8'd29;
        rom[228][9] = -8'd26;
        rom[228][10] = -8'd3;
        rom[228][11] = -8'd3;
        rom[228][12] = -8'd18;
        rom[228][13] = -8'd24;
        rom[228][14] = -8'd29;
        rom[228][15] = -8'd13;
        rom[228][16] = -8'd60;
        rom[228][17] = -8'd14;
        rom[228][18] = -8'd10;
        rom[228][19] = 8'd42;
        rom[228][20] = -8'd1;
        rom[228][21] = -8'd16;
        rom[228][22] = 8'd30;
        rom[228][23] = -8'd24;
        rom[228][24] = -8'd52;
        rom[228][25] = -8'd30;
        rom[228][26] = -8'd3;
        rom[228][27] = 8'd9;
        rom[228][28] = 8'd1;
        rom[228][29] = 8'd16;
        rom[228][30] = -8'd4;
        rom[228][31] = -8'd14;
        rom[228][32] = -8'd35;
        rom[228][33] = 8'd33;
        rom[228][34] = -8'd33;
        rom[228][35] = -8'd8;
        rom[228][36] = -8'd5;
        rom[228][37] = 8'd31;
        rom[228][38] = -8'd20;
        rom[228][39] = -8'd12;
        rom[228][40] = -8'd22;
        rom[228][41] = -8'd23;
        rom[228][42] = 8'd12;
        rom[228][43] = 8'd16;
        rom[228][44] = 8'd24;
        rom[228][45] = -8'd5;
        rom[228][46] = 8'd5;
        rom[228][47] = 8'd28;
        rom[228][48] = -8'd3;
        rom[228][49] = -8'd40;
        rom[228][50] = -8'd27;
        rom[228][51] = -8'd13;
        rom[228][52] = -8'd53;
        rom[228][53] = -8'd16;
        rom[228][54] = -8'd21;
        rom[228][55] = 8'd16;
        rom[228][56] = 8'd17;
        rom[228][57] = -8'd38;
        rom[228][58] = 8'd29;
        rom[228][59] = 8'd5;
        rom[228][60] = -8'd50;
        rom[228][61] = -8'd30;
        rom[228][62] = -8'd5;
        rom[228][63] = 8'd11;
        rom[229][0] = -8'd40;
        rom[229][1] = -8'd70;
        rom[229][2] = -8'd24;
        rom[229][3] = 8'd10;
        rom[229][4] = -8'd26;
        rom[229][5] = 8'd14;
        rom[229][6] = -8'd11;
        rom[229][7] = -8'd12;
        rom[229][8] = 8'd20;
        rom[229][9] = 8'd56;
        rom[229][10] = -8'd45;
        rom[229][11] = -8'd65;
        rom[229][12] = -8'd72;
        rom[229][13] = -8'd43;
        rom[229][14] = -8'd45;
        rom[229][15] = 8'd11;
        rom[229][16] = -8'd12;
        rom[229][17] = -8'd17;
        rom[229][18] = 8'd13;
        rom[229][19] = -8'd14;
        rom[229][20] = -8'd11;
        rom[229][21] = -8'd20;
        rom[229][22] = -8'd9;
        rom[229][23] = 8'd6;
        rom[229][24] = -8'd31;
        rom[229][25] = 8'd5;
        rom[229][26] = -8'd7;
        rom[229][27] = 8'd53;
        rom[229][28] = -8'd1;
        rom[229][29] = 8'd27;
        rom[229][30] = -8'd28;
        rom[229][31] = 8'd4;
        rom[229][32] = -8'd33;
        rom[229][33] = 8'd9;
        rom[229][34] = -8'd33;
        rom[229][35] = 8'd18;
        rom[229][36] = -8'd5;
        rom[229][37] = -8'd22;
        rom[229][38] = -8'd41;
        rom[229][39] = 8'd32;
        rom[229][40] = -8'd27;
        rom[229][41] = -8'd6;
        rom[229][42] = -8'd50;
        rom[229][43] = -8'd38;
        rom[229][44] = 8'd16;
        rom[229][45] = -8'd23;
        rom[229][46] = -8'd10;
        rom[229][47] = -8'd34;
        rom[229][48] = -8'd24;
        rom[229][49] = -8'd42;
        rom[229][50] = 8'd6;
        rom[229][51] = 8'd12;
        rom[229][52] = 8'd35;
        rom[229][53] = 8'd42;
        rom[229][54] = 8'd42;
        rom[229][55] = -8'd9;
        rom[229][56] = -8'd38;
        rom[229][57] = -8'd48;
        rom[229][58] = -8'd8;
        rom[229][59] = 8'd4;
        rom[229][60] = 8'd16;
        rom[229][61] = 8'd5;
        rom[229][62] = 8'd22;
        rom[229][63] = -8'd14;
        rom[230][0] = -8'd1;
        rom[230][1] = -8'd33;
        rom[230][2] = 8'd24;
        rom[230][3] = -8'd38;
        rom[230][4] = -8'd53;
        rom[230][5] = -8'd19;
        rom[230][6] = -8'd64;
        rom[230][7] = 8'd9;
        rom[230][8] = 8'd0;
        rom[230][9] = -8'd9;
        rom[230][10] = -8'd17;
        rom[230][11] = -8'd8;
        rom[230][12] = 8'd20;
        rom[230][13] = 8'd43;
        rom[230][14] = -8'd16;
        rom[230][15] = -8'd18;
        rom[230][16] = -8'd11;
        rom[230][17] = -8'd13;
        rom[230][18] = -8'd35;
        rom[230][19] = -8'd45;
        rom[230][20] = 8'd3;
        rom[230][21] = -8'd27;
        rom[230][22] = -8'd35;
        rom[230][23] = 8'd13;
        rom[230][24] = 8'd26;
        rom[230][25] = 8'd0;
        rom[230][26] = 8'd23;
        rom[230][27] = -8'd47;
        rom[230][28] = 8'd4;
        rom[230][29] = -8'd44;
        rom[230][30] = 8'd13;
        rom[230][31] = 8'd19;
        rom[230][32] = -8'd24;
        rom[230][33] = -8'd11;
        rom[230][34] = 8'd1;
        rom[230][35] = -8'd23;
        rom[230][36] = 8'd16;
        rom[230][37] = 8'd2;
        rom[230][38] = 8'd15;
        rom[230][39] = -8'd40;
        rom[230][40] = -8'd1;
        rom[230][41] = 8'd29;
        rom[230][42] = 8'd25;
        rom[230][43] = 8'd20;
        rom[230][44] = 8'd18;
        rom[230][45] = -8'd22;
        rom[230][46] = -8'd22;
        rom[230][47] = 8'd41;
        rom[230][48] = 8'd33;
        rom[230][49] = -8'd23;
        rom[230][50] = 8'd23;
        rom[230][51] = -8'd41;
        rom[230][52] = 8'd15;
        rom[230][53] = -8'd20;
        rom[230][54] = 8'd7;
        rom[230][55] = -8'd78;
        rom[230][56] = -8'd9;
        rom[230][57] = -8'd2;
        rom[230][58] = 8'd1;
        rom[230][59] = 8'd13;
        rom[230][60] = 8'd17;
        rom[230][61] = 8'd11;
        rom[230][62] = 8'd48;
        rom[230][63] = -8'd12;
        rom[231][0] = -8'd21;
        rom[231][1] = 8'd4;
        rom[231][2] = -8'd9;
        rom[231][3] = -8'd17;
        rom[231][4] = 8'd3;
        rom[231][5] = -8'd13;
        rom[231][6] = -8'd3;
        rom[231][7] = -8'd20;
        rom[231][8] = -8'd33;
        rom[231][9] = 8'd5;
        rom[231][10] = 8'd13;
        rom[231][11] = -8'd19;
        rom[231][12] = 8'd19;
        rom[231][13] = 8'd8;
        rom[231][14] = -8'd9;
        rom[231][15] = -8'd31;
        rom[231][16] = 8'd1;
        rom[231][17] = -8'd35;
        rom[231][18] = 8'd16;
        rom[231][19] = 8'd5;
        rom[231][20] = 8'd1;
        rom[231][21] = -8'd32;
        rom[231][22] = -8'd13;
        rom[231][23] = -8'd17;
        rom[231][24] = -8'd3;
        rom[231][25] = -8'd62;
        rom[231][26] = 8'd42;
        rom[231][27] = 8'd19;
        rom[231][28] = 8'd3;
        rom[231][29] = -8'd9;
        rom[231][30] = 8'd15;
        rom[231][31] = 8'd6;
        rom[231][32] = 8'd1;
        rom[231][33] = -8'd13;
        rom[231][34] = -8'd19;
        rom[231][35] = -8'd21;
        rom[231][36] = 8'd8;
        rom[231][37] = 8'd8;
        rom[231][38] = -8'd40;
        rom[231][39] = -8'd1;
        rom[231][40] = 8'd2;
        rom[231][41] = -8'd21;
        rom[231][42] = 8'd10;
        rom[231][43] = -8'd10;
        rom[231][44] = -8'd29;
        rom[231][45] = -8'd19;
        rom[231][46] = 8'd8;
        rom[231][47] = -8'd76;
        rom[231][48] = -8'd10;
        rom[231][49] = 8'd15;
        rom[231][50] = 8'd25;
        rom[231][51] = -8'd18;
        rom[231][52] = -8'd19;
        rom[231][53] = -8'd37;
        rom[231][54] = 8'd8;
        rom[231][55] = 8'd0;
        rom[231][56] = 8'd0;
        rom[231][57] = 8'd15;
        rom[231][58] = -8'd49;
        rom[231][59] = 8'd28;
        rom[231][60] = -8'd15;
        rom[231][61] = 8'd6;
        rom[231][62] = 8'd20;
        rom[231][63] = -8'd35;
        rom[232][0] = -8'd22;
        rom[232][1] = -8'd9;
        rom[232][2] = -8'd6;
        rom[232][3] = 8'd33;
        rom[232][4] = 8'd18;
        rom[232][5] = -8'd5;
        rom[232][6] = 8'd20;
        rom[232][7] = 8'd20;
        rom[232][8] = -8'd14;
        rom[232][9] = -8'd70;
        rom[232][10] = -8'd53;
        rom[232][11] = -8'd17;
        rom[232][12] = -8'd32;
        rom[232][13] = -8'd6;
        rom[232][14] = -8'd4;
        rom[232][15] = -8'd60;
        rom[232][16] = -8'd4;
        rom[232][17] = -8'd2;
        rom[232][18] = 8'd24;
        rom[232][19] = 8'd23;
        rom[232][20] = -8'd14;
        rom[232][21] = -8'd54;
        rom[232][22] = 8'd10;
        rom[232][23] = 8'd33;
        rom[232][24] = 8'd29;
        rom[232][25] = -8'd23;
        rom[232][26] = -8'd54;
        rom[232][27] = -8'd34;
        rom[232][28] = -8'd22;
        rom[232][29] = -8'd34;
        rom[232][30] = -8'd30;
        rom[232][31] = 8'd6;
        rom[232][32] = 8'd8;
        rom[232][33] = 8'd2;
        rom[232][34] = 8'd22;
        rom[232][35] = 8'd0;
        rom[232][36] = -8'd27;
        rom[232][37] = 8'd12;
        rom[232][38] = 8'd33;
        rom[232][39] = -8'd22;
        rom[232][40] = 8'd34;
        rom[232][41] = -8'd4;
        rom[232][42] = 8'd10;
        rom[232][43] = -8'd15;
        rom[232][44] = 8'd37;
        rom[232][45] = 8'd1;
        rom[232][46] = 8'd6;
        rom[232][47] = 8'd14;
        rom[232][48] = 8'd39;
        rom[232][49] = -8'd25;
        rom[232][50] = 8'd32;
        rom[232][51] = 8'd14;
        rom[232][52] = -8'd30;
        rom[232][53] = -8'd16;
        rom[232][54] = 8'd1;
        rom[232][55] = -8'd4;
        rom[232][56] = 8'd54;
        rom[232][57] = -8'd28;
        rom[232][58] = 8'd10;
        rom[232][59] = -8'd50;
        rom[232][60] = 8'd12;
        rom[232][61] = -8'd11;
        rom[232][62] = 8'd1;
        rom[232][63] = 8'd1;
        rom[233][0] = -8'd21;
        rom[233][1] = -8'd4;
        rom[233][2] = -8'd4;
        rom[233][3] = 8'd20;
        rom[233][4] = -8'd8;
        rom[233][5] = -8'd24;
        rom[233][6] = 8'd27;
        rom[233][7] = -8'd19;
        rom[233][8] = -8'd2;
        rom[233][9] = 8'd18;
        rom[233][10] = -8'd33;
        rom[233][11] = -8'd71;
        rom[233][12] = -8'd18;
        rom[233][13] = 8'd10;
        rom[233][14] = -8'd23;
        rom[233][15] = -8'd9;
        rom[233][16] = -8'd18;
        rom[233][17] = 8'd4;
        rom[233][18] = 8'd4;
        rom[233][19] = -8'd31;
        rom[233][20] = -8'd7;
        rom[233][21] = -8'd33;
        rom[233][22] = -8'd34;
        rom[233][23] = -8'd25;
        rom[233][24] = 8'd6;
        rom[233][25] = 8'd7;
        rom[233][26] = 8'd8;
        rom[233][27] = 8'd56;
        rom[233][28] = 8'd4;
        rom[233][29] = 8'd7;
        rom[233][30] = -8'd22;
        rom[233][31] = -8'd4;
        rom[233][32] = -8'd38;
        rom[233][33] = 8'd14;
        rom[233][34] = 8'd3;
        rom[233][35] = -8'd18;
        rom[233][36] = 8'd23;
        rom[233][37] = -8'd90;
        rom[233][38] = -8'd13;
        rom[233][39] = -8'd24;
        rom[233][40] = -8'd2;
        rom[233][41] = 8'd0;
        rom[233][42] = 8'd17;
        rom[233][43] = 8'd38;
        rom[233][44] = 8'd21;
        rom[233][45] = 8'd20;
        rom[233][46] = -8'd4;
        rom[233][47] = -8'd82;
        rom[233][48] = 8'd10;
        rom[233][49] = -8'd52;
        rom[233][50] = -8'd10;
        rom[233][51] = 8'd20;
        rom[233][52] = 8'd11;
        rom[233][53] = 8'd7;
        rom[233][54] = -8'd1;
        rom[233][55] = 8'd18;
        rom[233][56] = 8'd12;
        rom[233][57] = 8'd46;
        rom[233][58] = -8'd15;
        rom[233][59] = 8'd22;
        rom[233][60] = -8'd17;
        rom[233][61] = 8'd12;
        rom[233][62] = 8'd4;
        rom[233][63] = 8'd8;
        rom[234][0] = 8'd21;
        rom[234][1] = -8'd13;
        rom[234][2] = -8'd5;
        rom[234][3] = -8'd17;
        rom[234][4] = -8'd46;
        rom[234][5] = -8'd10;
        rom[234][6] = -8'd1;
        rom[234][7] = 8'd5;
        rom[234][8] = 8'd0;
        rom[234][9] = 8'd18;
        rom[234][10] = 8'd5;
        rom[234][11] = 8'd9;
        rom[234][12] = -8'd13;
        rom[234][13] = -8'd11;
        rom[234][14] = -8'd7;
        rom[234][15] = 8'd14;
        rom[234][16] = 8'd30;
        rom[234][17] = -8'd44;
        rom[234][18] = 8'd13;
        rom[234][19] = 8'd1;
        rom[234][20] = 8'd6;
        rom[234][21] = 8'd21;
        rom[234][22] = 8'd10;
        rom[234][23] = 8'd12;
        rom[234][24] = -8'd41;
        rom[234][25] = -8'd40;
        rom[234][26] = 8'd12;
        rom[234][27] = 8'd99;
        rom[234][28] = -8'd21;
        rom[234][29] = -8'd14;
        rom[234][30] = 8'd5;
        rom[234][31] = 8'd25;
        rom[234][32] = -8'd1;
        rom[234][33] = 8'd10;
        rom[234][34] = -8'd26;
        rom[234][35] = 8'd1;
        rom[234][36] = -8'd5;
        rom[234][37] = -8'd5;
        rom[234][38] = 8'd23;
        rom[234][39] = -8'd17;
        rom[234][40] = -8'd26;
        rom[234][41] = 8'd6;
        rom[234][42] = 8'd18;
        rom[234][43] = -8'd6;
        rom[234][44] = -8'd5;
        rom[234][45] = 8'd20;
        rom[234][46] = 8'd9;
        rom[234][47] = -8'd7;
        rom[234][48] = 8'd10;
        rom[234][49] = -8'd36;
        rom[234][50] = 8'd25;
        rom[234][51] = -8'd26;
        rom[234][52] = -8'd24;
        rom[234][53] = -8'd8;
        rom[234][54] = 8'd20;
        rom[234][55] = -8'd19;
        rom[234][56] = -8'd1;
        rom[234][57] = 8'd54;
        rom[234][58] = 8'd0;
        rom[234][59] = 8'd31;
        rom[234][60] = 8'd10;
        rom[234][61] = -8'd22;
        rom[234][62] = 8'd4;
        rom[234][63] = -8'd21;
        rom[235][0] = 8'd1;
        rom[235][1] = -8'd30;
        rom[235][2] = 8'd18;
        rom[235][3] = -8'd6;
        rom[235][4] = 8'd13;
        rom[235][5] = 8'd6;
        rom[235][6] = -8'd11;
        rom[235][7] = 8'd10;
        rom[235][8] = 8'd3;
        rom[235][9] = -8'd15;
        rom[235][10] = 8'd22;
        rom[235][11] = 8'd10;
        rom[235][12] = 8'd32;
        rom[235][13] = -8'd24;
        rom[235][14] = -8'd13;
        rom[235][15] = -8'd25;
        rom[235][16] = -8'd25;
        rom[235][17] = -8'd6;
        rom[235][18] = 8'd6;
        rom[235][19] = 8'd6;
        rom[235][20] = -8'd7;
        rom[235][21] = 8'd15;
        rom[235][22] = -8'd30;
        rom[235][23] = 8'd0;
        rom[235][24] = -8'd1;
        rom[235][25] = -8'd35;
        rom[235][26] = -8'd34;
        rom[235][27] = 8'd23;
        rom[235][28] = 8'd1;
        rom[235][29] = -8'd80;
        rom[235][30] = -8'd4;
        rom[235][31] = -8'd14;
        rom[235][32] = -8'd33;
        rom[235][33] = -8'd37;
        rom[235][34] = -8'd17;
        rom[235][35] = 8'd41;
        rom[235][36] = 8'd18;
        rom[235][37] = 8'd7;
        rom[235][38] = 8'd35;
        rom[235][39] = -8'd13;
        rom[235][40] = -8'd4;
        rom[235][41] = 8'd16;
        rom[235][42] = 8'd6;
        rom[235][43] = 8'd3;
        rom[235][44] = -8'd18;
        rom[235][45] = 8'd15;
        rom[235][46] = -8'd14;
        rom[235][47] = 8'd2;
        rom[235][48] = -8'd33;
        rom[235][49] = -8'd8;
        rom[235][50] = -8'd15;
        rom[235][51] = -8'd12;
        rom[235][52] = -8'd35;
        rom[235][53] = 8'd28;
        rom[235][54] = 8'd19;
        rom[235][55] = 8'd56;
        rom[235][56] = -8'd13;
        rom[235][57] = -8'd42;
        rom[235][58] = -8'd16;
        rom[235][59] = 8'd14;
        rom[235][60] = -8'd26;
        rom[235][61] = 8'd1;
        rom[235][62] = -8'd20;
        rom[235][63] = -8'd21;
        rom[236][0] = -8'd13;
        rom[236][1] = -8'd41;
        rom[236][2] = -8'd15;
        rom[236][3] = 8'd9;
        rom[236][4] = 8'd18;
        rom[236][5] = 8'd10;
        rom[236][6] = -8'd17;
        rom[236][7] = -8'd39;
        rom[236][8] = -8'd17;
        rom[236][9] = -8'd1;
        rom[236][10] = 8'd12;
        rom[236][11] = -8'd9;
        rom[236][12] = 8'd22;
        rom[236][13] = -8'd13;
        rom[236][14] = -8'd53;
        rom[236][15] = -8'd16;
        rom[236][16] = -8'd31;
        rom[236][17] = 8'd3;
        rom[236][18] = -8'd63;
        rom[236][19] = -8'd34;
        rom[236][20] = 8'd5;
        rom[236][21] = -8'd13;
        rom[236][22] = -8'd5;
        rom[236][23] = 8'd0;
        rom[236][24] = -8'd32;
        rom[236][25] = -8'd35;
        rom[236][26] = 8'd8;
        rom[236][27] = 8'd10;
        rom[236][28] = -8'd32;
        rom[236][29] = -8'd21;
        rom[236][30] = 8'd0;
        rom[236][31] = -8'd30;
        rom[236][32] = -8'd18;
        rom[236][33] = -8'd16;
        rom[236][34] = -8'd28;
        rom[236][35] = -8'd8;
        rom[236][36] = 8'd1;
        rom[236][37] = 8'd5;
        rom[236][38] = -8'd25;
        rom[236][39] = 8'd16;
        rom[236][40] = -8'd18;
        rom[236][41] = -8'd34;
        rom[236][42] = 8'd4;
        rom[236][43] = -8'd34;
        rom[236][44] = 8'd6;
        rom[236][45] = -8'd25;
        rom[236][46] = -8'd13;
        rom[236][47] = -8'd12;
        rom[236][48] = -8'd35;
        rom[236][49] = -8'd2;
        rom[236][50] = -8'd21;
        rom[236][51] = 8'd1;
        rom[236][52] = 8'd14;
        rom[236][53] = -8'd21;
        rom[236][54] = 8'd4;
        rom[236][55] = -8'd2;
        rom[236][56] = 8'd11;
        rom[236][57] = 8'd25;
        rom[236][58] = -8'd32;
        rom[236][59] = 8'd3;
        rom[236][60] = -8'd19;
        rom[236][61] = -8'd28;
        rom[236][62] = -8'd45;
        rom[236][63] = -8'd28;
        rom[237][0] = 8'd2;
        rom[237][1] = 8'd41;
        rom[237][2] = -8'd4;
        rom[237][3] = -8'd47;
        rom[237][4] = 8'd40;
        rom[237][5] = -8'd14;
        rom[237][6] = 8'd66;
        rom[237][7] = -8'd49;
        rom[237][8] = 8'd3;
        rom[237][9] = 8'd13;
        rom[237][10] = -8'd61;
        rom[237][11] = 8'd29;
        rom[237][12] = 8'd14;
        rom[237][13] = -8'd13;
        rom[237][14] = -8'd22;
        rom[237][15] = -8'd30;
        rom[237][16] = -8'd6;
        rom[237][17] = -8'd47;
        rom[237][18] = -8'd32;
        rom[237][19] = 8'd12;
        rom[237][20] = -8'd9;
        rom[237][21] = 8'd23;
        rom[237][22] = 8'd6;
        rom[237][23] = -8'd49;
        rom[237][24] = 8'd0;
        rom[237][25] = 8'd33;
        rom[237][26] = -8'd21;
        rom[237][27] = -8'd19;
        rom[237][28] = 8'd11;
        rom[237][29] = 8'd1;
        rom[237][30] = 8'd10;
        rom[237][31] = 8'd7;
        rom[237][32] = 8'd30;
        rom[237][33] = 8'd2;
        rom[237][34] = 8'd50;
        rom[237][35] = -8'd6;
        rom[237][36] = -8'd9;
        rom[237][37] = -8'd5;
        rom[237][38] = 8'd31;
        rom[237][39] = -8'd11;
        rom[237][40] = -8'd35;
        rom[237][41] = 8'd53;
        rom[237][42] = -8'd27;
        rom[237][43] = -8'd20;
        rom[237][44] = -8'd37;
        rom[237][45] = -8'd40;
        rom[237][46] = -8'd24;
        rom[237][47] = 8'd37;
        rom[237][48] = 8'd3;
        rom[237][49] = 8'd6;
        rom[237][50] = 8'd22;
        rom[237][51] = 8'd13;
        rom[237][52] = -8'd26;
        rom[237][53] = 8'd9;
        rom[237][54] = 8'd25;
        rom[237][55] = 8'd15;
        rom[237][56] = 8'd0;
        rom[237][57] = -8'd84;
        rom[237][58] = 8'd2;
        rom[237][59] = -8'd15;
        rom[237][60] = 8'd40;
        rom[237][61] = 8'd16;
        rom[237][62] = 8'd29;
        rom[237][63] = 8'd58;
        rom[238][0] = -8'd29;
        rom[238][1] = -8'd33;
        rom[238][2] = 8'd28;
        rom[238][3] = 8'd5;
        rom[238][4] = 8'd26;
        rom[238][5] = -8'd8;
        rom[238][6] = 8'd2;
        rom[238][7] = 8'd7;
        rom[238][8] = -8'd26;
        rom[238][9] = -8'd4;
        rom[238][10] = -8'd31;
        rom[238][11] = 8'd14;
        rom[238][12] = -8'd31;
        rom[238][13] = -8'd11;
        rom[238][14] = -8'd11;
        rom[238][15] = -8'd51;
        rom[238][16] = -8'd13;
        rom[238][17] = 8'd32;
        rom[238][18] = 8'd3;
        rom[238][19] = 8'd16;
        rom[238][20] = -8'd4;
        rom[238][21] = -8'd14;
        rom[238][22] = -8'd21;
        rom[238][23] = -8'd4;
        rom[238][24] = -8'd4;
        rom[238][25] = 8'd12;
        rom[238][26] = 8'd29;
        rom[238][27] = -8'd29;
        rom[238][28] = 8'd35;
        rom[238][29] = 8'd20;
        rom[238][30] = 8'd26;
        rom[238][31] = 8'd8;
        rom[238][32] = 8'd44;
        rom[238][33] = 8'd42;
        rom[238][34] = 8'd0;
        rom[238][35] = 8'd12;
        rom[238][36] = 8'd32;
        rom[238][37] = -8'd3;
        rom[238][38] = -8'd27;
        rom[238][39] = -8'd39;
        rom[238][40] = -8'd34;
        rom[238][41] = -8'd2;
        rom[238][42] = 8'd2;
        rom[238][43] = 8'd19;
        rom[238][44] = -8'd42;
        rom[238][45] = -8'd28;
        rom[238][46] = -8'd1;
        rom[238][47] = -8'd46;
        rom[238][48] = -8'd40;
        rom[238][49] = 8'd24;
        rom[238][50] = -8'd42;
        rom[238][51] = -8'd1;
        rom[238][52] = 8'd20;
        rom[238][53] = -8'd5;
        rom[238][54] = -8'd55;
        rom[238][55] = -8'd18;
        rom[238][56] = -8'd5;
        rom[238][57] = 8'd5;
        rom[238][58] = -8'd8;
        rom[238][59] = -8'd20;
        rom[238][60] = -8'd41;
        rom[238][61] = 8'd14;
        rom[238][62] = 8'd28;
        rom[238][63] = -8'd11;
        rom[239][0] = 8'd40;
        rom[239][1] = 8'd48;
        rom[239][2] = -8'd30;
        rom[239][3] = 8'd24;
        rom[239][4] = 8'd13;
        rom[239][5] = 8'd1;
        rom[239][6] = -8'd2;
        rom[239][7] = 8'd17;
        rom[239][8] = 8'd0;
        rom[239][9] = -8'd7;
        rom[239][10] = 8'd8;
        rom[239][11] = 8'd54;
        rom[239][12] = -8'd9;
        rom[239][13] = -8'd15;
        rom[239][14] = 8'd41;
        rom[239][15] = -8'd2;
        rom[239][16] = 8'd22;
        rom[239][17] = 8'd12;
        rom[239][18] = -8'd37;
        rom[239][19] = 8'd23;
        rom[239][20] = -8'd2;
        rom[239][21] = 8'd47;
        rom[239][22] = 8'd45;
        rom[239][23] = 8'd31;
        rom[239][24] = -8'd7;
        rom[239][25] = 8'd24;
        rom[239][26] = -8'd4;
        rom[239][27] = 8'd9;
        rom[239][28] = -8'd10;
        rom[239][29] = -8'd8;
        rom[239][30] = -8'd19;
        rom[239][31] = 8'd8;
        rom[239][32] = 8'd29;
        rom[239][33] = 8'd52;
        rom[239][34] = -8'd4;
        rom[239][35] = 8'd13;
        rom[239][36] = -8'd36;
        rom[239][37] = 8'd37;
        rom[239][38] = -8'd7;
        rom[239][39] = 8'd9;
        rom[239][40] = -8'd34;
        rom[239][41] = -8'd2;
        rom[239][42] = 8'd47;
        rom[239][43] = -8'd12;
        rom[239][44] = 8'd20;
        rom[239][45] = -8'd39;
        rom[239][46] = -8'd22;
        rom[239][47] = -8'd41;
        rom[239][48] = 8'd53;
        rom[239][49] = 8'd25;
        rom[239][50] = -8'd30;
        rom[239][51] = 8'd57;
        rom[239][52] = -8'd7;
        rom[239][53] = 8'd50;
        rom[239][54] = -8'd15;
        rom[239][55] = -8'd5;
        rom[239][56] = -8'd28;
        rom[239][57] = 8'd39;
        rom[239][58] = -8'd28;
        rom[239][59] = 8'd8;
        rom[239][60] = -8'd25;
        rom[239][61] = -8'd46;
        rom[239][62] = -8'd22;
        rom[239][63] = -8'd12;
        rom[240][0] = 8'd8;
        rom[240][1] = 8'd28;
        rom[240][2] = -8'd30;
        rom[240][3] = 8'd20;
        rom[240][4] = 8'd3;
        rom[240][5] = -8'd25;
        rom[240][6] = -8'd9;
        rom[240][7] = 8'd2;
        rom[240][8] = 8'd7;
        rom[240][9] = 8'd3;
        rom[240][10] = -8'd12;
        rom[240][11] = -8'd9;
        rom[240][12] = -8'd29;
        rom[240][13] = 8'd12;
        rom[240][14] = -8'd21;
        rom[240][15] = -8'd2;
        rom[240][16] = 8'd40;
        rom[240][17] = 8'd23;
        rom[240][18] = 8'd9;
        rom[240][19] = 8'd25;
        rom[240][20] = -8'd12;
        rom[240][21] = 8'd6;
        rom[240][22] = 8'd2;
        rom[240][23] = 8'd23;
        rom[240][24] = 8'd1;
        rom[240][25] = 8'd26;
        rom[240][26] = -8'd43;
        rom[240][27] = 8'd19;
        rom[240][28] = 8'd1;
        rom[240][29] = -8'd55;
        rom[240][30] = 8'd3;
        rom[240][31] = 8'd3;
        rom[240][32] = 8'd1;
        rom[240][33] = 8'd58;
        rom[240][34] = -8'd47;
        rom[240][35] = 8'd32;
        rom[240][36] = 8'd25;
        rom[240][37] = 8'd13;
        rom[240][38] = 8'd24;
        rom[240][39] = 8'd1;
        rom[240][40] = 8'd17;
        rom[240][41] = -8'd19;
        rom[240][42] = -8'd20;
        rom[240][43] = 8'd41;
        rom[240][44] = 8'd22;
        rom[240][45] = 8'd66;
        rom[240][46] = 8'd12;
        rom[240][47] = 8'd3;
        rom[240][48] = -8'd35;
        rom[240][49] = -8'd22;
        rom[240][50] = 8'd17;
        rom[240][51] = -8'd1;
        rom[240][52] = -8'd68;
        rom[240][53] = -8'd23;
        rom[240][54] = -8'd13;
        rom[240][55] = -8'd1;
        rom[240][56] = 8'd5;
        rom[240][57] = -8'd27;
        rom[240][58] = -8'd33;
        rom[240][59] = 8'd22;
        rom[240][60] = -8'd42;
        rom[240][61] = -8'd2;
        rom[240][62] = -8'd3;
        rom[240][63] = -8'd16;
        rom[241][0] = -8'd16;
        rom[241][1] = -8'd54;
        rom[241][2] = 8'd20;
        rom[241][3] = -8'd19;
        rom[241][4] = 8'd13;
        rom[241][5] = -8'd26;
        rom[241][6] = -8'd64;
        rom[241][7] = -8'd21;
        rom[241][8] = -8'd4;
        rom[241][9] = 8'd31;
        rom[241][10] = -8'd4;
        rom[241][11] = 8'd21;
        rom[241][12] = 8'd44;
        rom[241][13] = 8'd23;
        rom[241][14] = -8'd9;
        rom[241][15] = 8'd32;
        rom[241][16] = -8'd11;
        rom[241][17] = -8'd20;
        rom[241][18] = -8'd37;
        rom[241][19] = 8'd14;
        rom[241][20] = -8'd4;
        rom[241][21] = -8'd20;
        rom[241][22] = 8'd12;
        rom[241][23] = 8'd11;
        rom[241][24] = -8'd4;
        rom[241][25] = -8'd32;
        rom[241][26] = -8'd36;
        rom[241][27] = -8'd36;
        rom[241][28] = -8'd2;
        rom[241][29] = -8'd9;
        rom[241][30] = 8'd23;
        rom[241][31] = -8'd11;
        rom[241][32] = 8'd13;
        rom[241][33] = 8'd33;
        rom[241][34] = 8'd25;
        rom[241][35] = -8'd32;
        rom[241][36] = -8'd12;
        rom[241][37] = -8'd26;
        rom[241][38] = -8'd2;
        rom[241][39] = -8'd23;
        rom[241][40] = -8'd4;
        rom[241][41] = 8'd23;
        rom[241][42] = 8'd38;
        rom[241][43] = 8'd18;
        rom[241][44] = 8'd27;
        rom[241][45] = 8'd42;
        rom[241][46] = -8'd26;
        rom[241][47] = -8'd4;
        rom[241][48] = -8'd2;
        rom[241][49] = 8'd20;
        rom[241][50] = 8'd0;
        rom[241][51] = -8'd27;
        rom[241][52] = -8'd1;
        rom[241][53] = 8'd12;
        rom[241][54] = 8'd12;
        rom[241][55] = -8'd17;
        rom[241][56] = 8'd23;
        rom[241][57] = 8'd12;
        rom[241][58] = 8'd12;
        rom[241][59] = 8'd24;
        rom[241][60] = -8'd25;
        rom[241][61] = -8'd18;
        rom[241][62] = -8'd16;
        rom[241][63] = 8'd7;
        rom[242][0] = -8'd9;
        rom[242][1] = 8'd25;
        rom[242][2] = 8'd0;
        rom[242][3] = -8'd17;
        rom[242][4] = -8'd6;
        rom[242][5] = 8'd4;
        rom[242][6] = 8'd4;
        rom[242][7] = 8'd10;
        rom[242][8] = -8'd51;
        rom[242][9] = 8'd15;
        rom[242][10] = -8'd28;
        rom[242][11] = -8'd29;
        rom[242][12] = 8'd38;
        rom[242][13] = -8'd5;
        rom[242][14] = -8'd31;
        rom[242][15] = -8'd21;
        rom[242][16] = -8'd48;
        rom[242][17] = -8'd9;
        rom[242][18] = 8'd12;
        rom[242][19] = 8'd1;
        rom[242][20] = -8'd1;
        rom[242][21] = 8'd13;
        rom[242][22] = 8'd16;
        rom[242][23] = -8'd11;
        rom[242][24] = 8'd17;
        rom[242][25] = -8'd8;
        rom[242][26] = 8'd22;
        rom[242][27] = -8'd13;
        rom[242][28] = 8'd28;
        rom[242][29] = 8'd51;
        rom[242][30] = -8'd1;
        rom[242][31] = -8'd64;
        rom[242][32] = 8'd8;
        rom[242][33] = -8'd37;
        rom[242][34] = 8'd37;
        rom[242][35] = 8'd0;
        rom[242][36] = 8'd16;
        rom[242][37] = 8'd7;
        rom[242][38] = -8'd37;
        rom[242][39] = -8'd45;
        rom[242][40] = -8'd16;
        rom[242][41] = -8'd21;
        rom[242][42] = -8'd4;
        rom[242][43] = 8'd6;
        rom[242][44] = 8'd2;
        rom[242][45] = -8'd28;
        rom[242][46] = -8'd25;
        rom[242][47] = -8'd1;
        rom[242][48] = -8'd41;
        rom[242][49] = 8'd8;
        rom[242][50] = -8'd34;
        rom[242][51] = -8'd48;
        rom[242][52] = 8'd32;
        rom[242][53] = -8'd10;
        rom[242][54] = -8'd11;
        rom[242][55] = -8'd35;
        rom[242][56] = 8'd2;
        rom[242][57] = -8'd14;
        rom[242][58] = 8'd3;
        rom[242][59] = -8'd26;
        rom[242][60] = 8'd3;
        rom[242][61] = -8'd1;
        rom[242][62] = 8'd19;
        rom[242][63] = 8'd4;
        rom[243][0] = 8'd13;
        rom[243][1] = -8'd57;
        rom[243][2] = 8'd21;
        rom[243][3] = -8'd24;
        rom[243][4] = -8'd8;
        rom[243][5] = 8'd0;
        rom[243][6] = 8'd11;
        rom[243][7] = 8'd0;
        rom[243][8] = -8'd23;
        rom[243][9] = 8'd10;
        rom[243][10] = -8'd8;
        rom[243][11] = -8'd31;
        rom[243][12] = 8'd14;
        rom[243][13] = -8'd33;
        rom[243][14] = -8'd11;
        rom[243][15] = 8'd39;
        rom[243][16] = -8'd10;
        rom[243][17] = -8'd3;
        rom[243][18] = -8'd19;
        rom[243][19] = 8'd4;
        rom[243][20] = 8'd2;
        rom[243][21] = -8'd8;
        rom[243][22] = -8'd18;
        rom[243][23] = -8'd17;
        rom[243][24] = 8'd10;
        rom[243][25] = 8'd19;
        rom[243][26] = 8'd0;
        rom[243][27] = -8'd20;
        rom[243][28] = 8'd13;
        rom[243][29] = 8'd14;
        rom[243][30] = -8'd51;
        rom[243][31] = 8'd18;
        rom[243][32] = -8'd15;
        rom[243][33] = -8'd39;
        rom[243][34] = 8'd2;
        rom[243][35] = -8'd24;
        rom[243][36] = 8'd15;
        rom[243][37] = 8'd14;
        rom[243][38] = -8'd31;
        rom[243][39] = -8'd3;
        rom[243][40] = -8'd40;
        rom[243][41] = -8'd2;
        rom[243][42] = -8'd23;
        rom[243][43] = -8'd50;
        rom[243][44] = 8'd10;
        rom[243][45] = -8'd64;
        rom[243][46] = -8'd14;
        rom[243][47] = -8'd38;
        rom[243][48] = 8'd8;
        rom[243][49] = -8'd11;
        rom[243][50] = -8'd32;
        rom[243][51] = -8'd31;
        rom[243][52] = 8'd24;
        rom[243][53] = -8'd11;
        rom[243][54] = -8'd23;
        rom[243][55] = -8'd15;
        rom[243][56] = -8'd40;
        rom[243][57] = 8'd25;
        rom[243][58] = 8'd6;
        rom[243][59] = 8'd19;
        rom[243][60] = 8'd6;
        rom[243][61] = -8'd19;
        rom[243][62] = 8'd29;
        rom[243][63] = 8'd41;
        rom[244][0] = 8'd34;
        rom[244][1] = -8'd99;
        rom[244][2] = -8'd45;
        rom[244][3] = -8'd18;
        rom[244][4] = -8'd7;
        rom[244][5] = -8'd25;
        rom[244][6] = -8'd75;
        rom[244][7] = -8'd22;
        rom[244][8] = -8'd51;
        rom[244][9] = -8'd45;
        rom[244][10] = 8'd2;
        rom[244][11] = 8'd14;
        rom[244][12] = -8'd61;
        rom[244][13] = 8'd18;
        rom[244][14] = 8'd26;
        rom[244][15] = -8'd43;
        rom[244][16] = -8'd57;
        rom[244][17] = 8'd14;
        rom[244][18] = -8'd15;
        rom[244][19] = 8'd13;
        rom[244][20] = -8'd9;
        rom[244][21] = -8'd43;
        rom[244][22] = -8'd51;
        rom[244][23] = -8'd13;
        rom[244][24] = -8'd29;
        rom[244][25] = 8'd21;
        rom[244][26] = 8'd12;
        rom[244][27] = -8'd56;
        rom[244][28] = -8'd20;
        rom[244][29] = -8'd45;
        rom[244][30] = -8'd33;
        rom[244][31] = 8'd13;
        rom[244][32] = -8'd5;
        rom[244][33] = 8'd7;
        rom[244][34] = 8'd5;
        rom[244][35] = -8'd9;
        rom[244][36] = -8'd38;
        rom[244][37] = -8'd11;
        rom[244][38] = -8'd54;
        rom[244][39] = 8'd7;
        rom[244][40] = -8'd20;
        rom[244][41] = 8'd10;
        rom[244][42] = -8'd54;
        rom[244][43] = -8'd26;
        rom[244][44] = 8'd14;
        rom[244][45] = 8'd5;
        rom[244][46] = -8'd1;
        rom[244][47] = 8'd5;
        rom[244][48] = -8'd25;
        rom[244][49] = 8'd30;
        rom[244][50] = -8'd19;
        rom[244][51] = 8'd24;
        rom[244][52] = 8'd28;
        rom[244][53] = -8'd13;
        rom[244][54] = -8'd64;
        rom[244][55] = 8'd4;
        rom[244][56] = -8'd24;
        rom[244][57] = 8'd22;
        rom[244][58] = -8'd3;
        rom[244][59] = -8'd65;
        rom[244][60] = -8'd17;
        rom[244][61] = -8'd23;
        rom[244][62] = -8'd25;
        rom[244][63] = -8'd48;
        rom[245][0] = 8'd19;
        rom[245][1] = 8'd4;
        rom[245][2] = 8'd22;
        rom[245][3] = -8'd29;
        rom[245][4] = -8'd12;
        rom[245][5] = 8'd19;
        rom[245][6] = -8'd23;
        rom[245][7] = 8'd7;
        rom[245][8] = -8'd22;
        rom[245][9] = -8'd19;
        rom[245][10] = -8'd45;
        rom[245][11] = -8'd22;
        rom[245][12] = -8'd17;
        rom[245][13] = 8'd2;
        rom[245][14] = 8'd55;
        rom[245][15] = 8'd21;
        rom[245][16] = 8'd23;
        rom[245][17] = 8'd12;
        rom[245][18] = 8'd27;
        rom[245][19] = 8'd19;
        rom[245][20] = -8'd10;
        rom[245][21] = -8'd5;
        rom[245][22] = 8'd2;
        rom[245][23] = 8'd8;
        rom[245][24] = -8'd28;
        rom[245][25] = -8'd7;
        rom[245][26] = -8'd15;
        rom[245][27] = -8'd1;
        rom[245][28] = -8'd37;
        rom[245][29] = 8'd19;
        rom[245][30] = 8'd34;
        rom[245][31] = 8'd11;
        rom[245][32] = -8'd42;
        rom[245][33] = -8'd4;
        rom[245][34] = -8'd47;
        rom[245][35] = -8'd22;
        rom[245][36] = -8'd11;
        rom[245][37] = 8'd13;
        rom[245][38] = 8'd33;
        rom[245][39] = -8'd30;
        rom[245][40] = -8'd33;
        rom[245][41] = -8'd13;
        rom[245][42] = 8'd4;
        rom[245][43] = -8'd57;
        rom[245][44] = -8'd29;
        rom[245][45] = 8'd24;
        rom[245][46] = -8'd2;
        rom[245][47] = 8'd19;
        rom[245][48] = 8'd1;
        rom[245][49] = -8'd62;
        rom[245][50] = 8'd11;
        rom[245][51] = 8'd11;
        rom[245][52] = -8'd16;
        rom[245][53] = -8'd24;
        rom[245][54] = -8'd16;
        rom[245][55] = 8'd11;
        rom[245][56] = -8'd14;
        rom[245][57] = -8'd6;
        rom[245][58] = -8'd7;
        rom[245][59] = 8'd24;
        rom[245][60] = 8'd3;
        rom[245][61] = 8'd30;
        rom[245][62] = -8'd1;
        rom[245][63] = -8'd12;
        rom[246][0] = -8'd6;
        rom[246][1] = -8'd6;
        rom[246][2] = 8'd2;
        rom[246][3] = 8'd0;
        rom[246][4] = -8'd9;
        rom[246][5] = 8'd10;
        rom[246][6] = 8'd1;
        rom[246][7] = -8'd11;
        rom[246][8] = 8'd8;
        rom[246][9] = -8'd5;
        rom[246][10] = -8'd2;
        rom[246][11] = 8'd5;
        rom[246][12] = 8'd5;
        rom[246][13] = -8'd9;
        rom[246][14] = 8'd13;
        rom[246][15] = -8'd3;
        rom[246][16] = 8'd8;
        rom[246][17] = -8'd4;
        rom[246][18] = -8'd7;
        rom[246][19] = 8'd12;
        rom[246][20] = -8'd3;
        rom[246][21] = -8'd6;
        rom[246][22] = 8'd6;
        rom[246][23] = 8'd7;
        rom[246][24] = -8'd8;
        rom[246][25] = -8'd16;
        rom[246][26] = -8'd15;
        rom[246][27] = -8'd5;
        rom[246][28] = 8'd3;
        rom[246][29] = 8'd5;
        rom[246][30] = 8'd5;
        rom[246][31] = -8'd7;
        rom[246][32] = -8'd14;
        rom[246][33] = -8'd11;
        rom[246][34] = -8'd2;
        rom[246][35] = 8'd7;
        rom[246][36] = -8'd3;
        rom[246][37] = 8'd5;
        rom[246][38] = 8'd1;
        rom[246][39] = 8'd8;
        rom[246][40] = 8'd8;
        rom[246][41] = -8'd7;
        rom[246][42] = -8'd1;
        rom[246][43] = -8'd1;
        rom[246][44] = -8'd7;
        rom[246][45] = 8'd4;
        rom[246][46] = -8'd4;
        rom[246][47] = 8'd0;
        rom[246][48] = 8'd0;
        rom[246][49] = -8'd7;
        rom[246][50] = -8'd1;
        rom[246][51] = 8'd6;
        rom[246][52] = 8'd3;
        rom[246][53] = -8'd3;
        rom[246][54] = -8'd2;
        rom[246][55] = -8'd6;
        rom[246][56] = -8'd7;
        rom[246][57] = 8'd5;
        rom[246][58] = 8'd1;
        rom[246][59] = -8'd3;
        rom[246][60] = 8'd2;
        rom[246][61] = 8'd6;
        rom[246][62] = 8'd9;
        rom[246][63] = -8'd7;
        rom[247][0] = 8'd47;
        rom[247][1] = 8'd9;
        rom[247][2] = -8'd4;
        rom[247][3] = 8'd10;
        rom[247][4] = 8'd40;
        rom[247][5] = -8'd18;
        rom[247][6] = -8'd15;
        rom[247][7] = -8'd25;
        rom[247][8] = 8'd24;
        rom[247][9] = 8'd6;
        rom[247][10] = -8'd3;
        rom[247][11] = -8'd8;
        rom[247][12] = 8'd1;
        rom[247][13] = 8'd2;
        rom[247][14] = -8'd5;
        rom[247][15] = -8'd16;
        rom[247][16] = -8'd11;
        rom[247][17] = 8'd15;
        rom[247][18] = -8'd32;
        rom[247][19] = -8'd42;
        rom[247][20] = -8'd1;
        rom[247][21] = -8'd13;
        rom[247][22] = 8'd45;
        rom[247][23] = 8'd10;
        rom[247][24] = -8'd64;
        rom[247][25] = 8'd10;
        rom[247][26] = -8'd14;
        rom[247][27] = -8'd42;
        rom[247][28] = -8'd20;
        rom[247][29] = 8'd8;
        rom[247][30] = -8'd36;
        rom[247][31] = 8'd8;
        rom[247][32] = -8'd3;
        rom[247][33] = 8'd3;
        rom[247][34] = 8'd23;
        rom[247][35] = -8'd39;
        rom[247][36] = -8'd28;
        rom[247][37] = 8'd23;
        rom[247][38] = -8'd42;
        rom[247][39] = -8'd9;
        rom[247][40] = 8'd29;
        rom[247][41] = 8'd17;
        rom[247][42] = -8'd30;
        rom[247][43] = -8'd35;
        rom[247][44] = 8'd22;
        rom[247][45] = -8'd11;
        rom[247][46] = 8'd7;
        rom[247][47] = 8'd2;
        rom[247][48] = 8'd0;
        rom[247][49] = 8'd20;
        rom[247][50] = -8'd4;
        rom[247][51] = 8'd2;
        rom[247][52] = 8'd7;
        rom[247][53] = -8'd5;
        rom[247][54] = -8'd11;
        rom[247][55] = -8'd45;
        rom[247][56] = 8'd6;
        rom[247][57] = 8'd4;
        rom[247][58] = 8'd17;
        rom[247][59] = 8'd1;
        rom[247][60] = -8'd66;
        rom[247][61] = 8'd6;
        rom[247][62] = 8'd14;
        rom[247][63] = 8'd20;
        rom[248][0] = 8'd17;
        rom[248][1] = 8'd28;
        rom[248][2] = -8'd9;
        rom[248][3] = -8'd32;
        rom[248][4] = -8'd15;
        rom[248][5] = -8'd1;
        rom[248][6] = 8'd4;
        rom[248][7] = -8'd2;
        rom[248][8] = 8'd5;
        rom[248][9] = -8'd26;
        rom[248][10] = 8'd18;
        rom[248][11] = 8'd2;
        rom[248][12] = 8'd0;
        rom[248][13] = 8'd5;
        rom[248][14] = -8'd16;
        rom[248][15] = 8'd25;
        rom[248][16] = 8'd24;
        rom[248][17] = -8'd21;
        rom[248][18] = 8'd11;
        rom[248][19] = -8'd26;
        rom[248][20] = -8'd6;
        rom[248][21] = 8'd7;
        rom[248][22] = 8'd21;
        rom[248][23] = 8'd26;
        rom[248][24] = -8'd45;
        rom[248][25] = 8'd3;
        rom[248][26] = 8'd23;
        rom[248][27] = -8'd14;
        rom[248][28] = -8'd23;
        rom[248][29] = 8'd7;
        rom[248][30] = 8'd1;
        rom[248][31] = -8'd7;
        rom[248][32] = -8'd16;
        rom[248][33] = -8'd58;
        rom[248][34] = 8'd9;
        rom[248][35] = -8'd4;
        rom[248][36] = -8'd9;
        rom[248][37] = -8'd2;
        rom[248][38] = -8'd9;
        rom[248][39] = -8'd8;
        rom[248][40] = 8'd7;
        rom[248][41] = -8'd20;
        rom[248][42] = -8'd42;
        rom[248][43] = -8'd27;
        rom[248][44] = -8'd2;
        rom[248][45] = -8'd27;
        rom[248][46] = -8'd10;
        rom[248][47] = 8'd11;
        rom[248][48] = -8'd18;
        rom[248][49] = 8'd8;
        rom[248][50] = -8'd31;
        rom[248][51] = 8'd9;
        rom[248][52] = 8'd12;
        rom[248][53] = -8'd3;
        rom[248][54] = 8'd13;
        rom[248][55] = -8'd10;
        rom[248][56] = 8'd15;
        rom[248][57] = -8'd3;
        rom[248][58] = -8'd43;
        rom[248][59] = 8'd8;
        rom[248][60] = 8'd11;
        rom[248][61] = 8'd9;
        rom[248][62] = 8'd19;
        rom[248][63] = 8'd1;
        rom[249][0] = 8'd38;
        rom[249][1] = -8'd2;
        rom[249][2] = 8'd15;
        rom[249][3] = 8'd18;
        rom[249][4] = -8'd5;
        rom[249][5] = 8'd22;
        rom[249][6] = 8'd40;
        rom[249][7] = 8'd11;
        rom[249][8] = -8'd10;
        rom[249][9] = -8'd17;
        rom[249][10] = 8'd9;
        rom[249][11] = -8'd34;
        rom[249][12] = 8'd10;
        rom[249][13] = 8'd3;
        rom[249][14] = -8'd38;
        rom[249][15] = 8'd10;
        rom[249][16] = -8'd10;
        rom[249][17] = -8'd15;
        rom[249][18] = -8'd2;
        rom[249][19] = 8'd4;
        rom[249][20] = -8'd12;
        rom[249][21] = 8'd14;
        rom[249][22] = -8'd25;
        rom[249][23] = 8'd15;
        rom[249][24] = 8'd3;
        rom[249][25] = -8'd3;
        rom[249][26] = 8'd34;
        rom[249][27] = -8'd5;
        rom[249][28] = 8'd16;
        rom[249][29] = 8'd21;
        rom[249][30] = -8'd24;
        rom[249][31] = 8'd34;
        rom[249][32] = 8'd1;
        rom[249][33] = -8'd4;
        rom[249][34] = 8'd14;
        rom[249][35] = -8'd14;
        rom[249][36] = 8'd20;
        rom[249][37] = 8'd29;
        rom[249][38] = 8'd5;
        rom[249][39] = -8'd6;
        rom[249][40] = -8'd30;
        rom[249][41] = -8'd52;
        rom[249][42] = 8'd14;
        rom[249][43] = 8'd5;
        rom[249][44] = -8'd19;
        rom[249][45] = -8'd21;
        rom[249][46] = 8'd19;
        rom[249][47] = 8'd45;
        rom[249][48] = -8'd55;
        rom[249][49] = -8'd12;
        rom[249][50] = 8'd7;
        rom[249][51] = -8'd23;
        rom[249][52] = 8'd19;
        rom[249][53] = -8'd46;
        rom[249][54] = -8'd26;
        rom[249][55] = 8'd2;
        rom[249][56] = -8'd26;
        rom[249][57] = 8'd58;
        rom[249][58] = 8'd21;
        rom[249][59] = 8'd10;
        rom[249][60] = 8'd17;
        rom[249][61] = -8'd20;
        rom[249][62] = 8'd39;
        rom[249][63] = -8'd3;
        rom[250][0] = -8'd5;
        rom[250][1] = 8'd24;
        rom[250][2] = 8'd4;
        rom[250][3] = 8'd30;
        rom[250][4] = -8'd23;
        rom[250][5] = -8'd26;
        rom[250][6] = -8'd24;
        rom[250][7] = 8'd15;
        rom[250][8] = -8'd2;
        rom[250][9] = -8'd1;
        rom[250][10] = 8'd35;
        rom[250][11] = -8'd16;
        rom[250][12] = 8'd7;
        rom[250][13] = 8'd9;
        rom[250][14] = -8'd23;
        rom[250][15] = 8'd43;
        rom[250][16] = 8'd5;
        rom[250][17] = 8'd31;
        rom[250][18] = -8'd34;
        rom[250][19] = -8'd9;
        rom[250][20] = -8'd15;
        rom[250][21] = -8'd10;
        rom[250][22] = 8'd6;
        rom[250][23] = 8'd13;
        rom[250][24] = -8'd9;
        rom[250][25] = 8'd8;
        rom[250][26] = 8'd4;
        rom[250][27] = -8'd17;
        rom[250][28] = 8'd40;
        rom[250][29] = -8'd7;
        rom[250][30] = 8'd10;
        rom[250][31] = -8'd7;
        rom[250][32] = 8'd26;
        rom[250][33] = -8'd13;
        rom[250][34] = 8'd17;
        rom[250][35] = -8'd35;
        rom[250][36] = -8'd1;
        rom[250][37] = 8'd35;
        rom[250][38] = -8'd42;
        rom[250][39] = -8'd54;
        rom[250][40] = -8'd6;
        rom[250][41] = -8'd13;
        rom[250][42] = -8'd10;
        rom[250][43] = 8'd38;
        rom[250][44] = -8'd3;
        rom[250][45] = -8'd61;
        rom[250][46] = 8'd3;
        rom[250][47] = 8'd0;
        rom[250][48] = -8'd38;
        rom[250][49] = 8'd0;
        rom[250][50] = -8'd65;
        rom[250][51] = -8'd85;
        rom[250][52] = 8'd54;
        rom[250][53] = -8'd4;
        rom[250][54] = -8'd16;
        rom[250][55] = -8'd19;
        rom[250][56] = 8'd13;
        rom[250][57] = 8'd2;
        rom[250][58] = 8'd1;
        rom[250][59] = -8'd13;
        rom[250][60] = 8'd21;
        rom[250][61] = -8'd13;
        rom[250][62] = -8'd24;
        rom[250][63] = -8'd38;
        rom[251][0] = -8'd8;
        rom[251][1] = 8'd15;
        rom[251][2] = -8'd13;
        rom[251][3] = -8'd16;
        rom[251][4] = -8'd20;
        rom[251][5] = 8'd15;
        rom[251][6] = -8'd35;
        rom[251][7] = 8'd1;
        rom[251][8] = -8'd13;
        rom[251][9] = 8'd5;
        rom[251][10] = 8'd25;
        rom[251][11] = 8'd12;
        rom[251][12] = 8'd8;
        rom[251][13] = 8'd8;
        rom[251][14] = 8'd17;
        rom[251][15] = -8'd60;
        rom[251][16] = 8'd11;
        rom[251][17] = 8'd2;
        rom[251][18] = 8'd2;
        rom[251][19] = -8'd10;
        rom[251][20] = 8'd1;
        rom[251][21] = -8'd29;
        rom[251][22] = 8'd10;
        rom[251][23] = 8'd20;
        rom[251][24] = -8'd38;
        rom[251][25] = -8'd49;
        rom[251][26] = -8'd22;
        rom[251][27] = -8'd8;
        rom[251][28] = -8'd13;
        rom[251][29] = -8'd61;
        rom[251][30] = -8'd25;
        rom[251][31] = -8'd42;
        rom[251][32] = -8'd65;
        rom[251][33] = -8'd8;
        rom[251][34] = -8'd10;
        rom[251][35] = 8'd1;
        rom[251][36] = -8'd10;
        rom[251][37] = 8'd27;
        rom[251][38] = -8'd5;
        rom[251][39] = -8'd1;
        rom[251][40] = 8'd1;
        rom[251][41] = -8'd20;
        rom[251][42] = -8'd19;
        rom[251][43] = 8'd16;
        rom[251][44] = 8'd1;
        rom[251][45] = 8'd3;
        rom[251][46] = -8'd46;
        rom[251][47] = 8'd7;
        rom[251][48] = -8'd16;
        rom[251][49] = -8'd5;
        rom[251][50] = -8'd55;
        rom[251][51] = -8'd22;
        rom[251][52] = -8'd8;
        rom[251][53] = 8'd6;
        rom[251][54] = -8'd23;
        rom[251][55] = -8'd8;
        rom[251][56] = -8'd25;
        rom[251][57] = -8'd74;
        rom[251][58] = 8'd15;
        rom[251][59] = -8'd15;
        rom[251][60] = 8'd25;
        rom[251][61] = -8'd52;
        rom[251][62] = -8'd19;
        rom[251][63] = -8'd15;
        rom[252][0] = -8'd9;
        rom[252][1] = 8'd8;
        rom[252][2] = -8'd26;
        rom[252][3] = 8'd21;
        rom[252][4] = 8'd25;
        rom[252][5] = -8'd55;
        rom[252][6] = 8'd4;
        rom[252][7] = -8'd18;
        rom[252][8] = 8'd18;
        rom[252][9] = -8'd18;
        rom[252][10] = -8'd33;
        rom[252][11] = -8'd8;
        rom[252][12] = 8'd10;
        rom[252][13] = -8'd47;
        rom[252][14] = -8'd30;
        rom[252][15] = 8'd13;
        rom[252][16] = -8'd34;
        rom[252][17] = -8'd1;
        rom[252][18] = -8'd19;
        rom[252][19] = -8'd1;
        rom[252][20] = -8'd11;
        rom[252][21] = -8'd31;
        rom[252][22] = -8'd24;
        rom[252][23] = 8'd23;
        rom[252][24] = -8'd28;
        rom[252][25] = 8'd9;
        rom[252][26] = 8'd16;
        rom[252][27] = 8'd30;
        rom[252][28] = 8'd16;
        rom[252][29] = 8'd3;
        rom[252][30] = 8'd2;
        rom[252][31] = 8'd5;
        rom[252][32] = -8'd2;
        rom[252][33] = -8'd25;
        rom[252][34] = 8'd29;
        rom[252][35] = -8'd14;
        rom[252][36] = -8'd14;
        rom[252][37] = 8'd27;
        rom[252][38] = -8'd11;
        rom[252][39] = -8'd8;
        rom[252][40] = -8'd23;
        rom[252][41] = -8'd10;
        rom[252][42] = -8'd55;
        rom[252][43] = 8'd27;
        rom[252][44] = 8'd25;
        rom[252][45] = -8'd26;
        rom[252][46] = -8'd2;
        rom[252][47] = -8'd34;
        rom[252][48] = -8'd59;
        rom[252][49] = -8'd29;
        rom[252][50] = 8'd18;
        rom[252][51] = -8'd11;
        rom[252][52] = 8'd2;
        rom[252][53] = -8'd17;
        rom[252][54] = 8'd11;
        rom[252][55] = -8'd33;
        rom[252][56] = 8'd0;
        rom[252][57] = -8'd30;
        rom[252][58] = -8'd25;
        rom[252][59] = -8'd33;
        rom[252][60] = -8'd19;
        rom[252][61] = -8'd71;
        rom[252][62] = 8'd32;
        rom[252][63] = -8'd15;
        rom[253][0] = 8'd4;
        rom[253][1] = -8'd23;
        rom[253][2] = 8'd6;
        rom[253][3] = -8'd46;
        rom[253][4] = 8'd10;
        rom[253][5] = 8'd21;
        rom[253][6] = -8'd49;
        rom[253][7] = -8'd12;
        rom[253][8] = -8'd20;
        rom[253][9] = -8'd27;
        rom[253][10] = 8'd21;
        rom[253][11] = 8'd12;
        rom[253][12] = -8'd17;
        rom[253][13] = 8'd25;
        rom[253][14] = -8'd29;
        rom[253][15] = -8'd7;
        rom[253][16] = 8'd2;
        rom[253][17] = -8'd23;
        rom[253][18] = 8'd11;
        rom[253][19] = -8'd7;
        rom[253][20] = -8'd11;
        rom[253][21] = 8'd18;
        rom[253][22] = -8'd1;
        rom[253][23] = 8'd6;
        rom[253][24] = -8'd14;
        rom[253][25] = -8'd39;
        rom[253][26] = 8'd33;
        rom[253][27] = -8'd50;
        rom[253][28] = -8'd7;
        rom[253][29] = -8'd7;
        rom[253][30] = 8'd20;
        rom[253][31] = 8'd3;
        rom[253][32] = 8'd13;
        rom[253][33] = -8'd1;
        rom[253][34] = 8'd16;
        rom[253][35] = 8'd28;
        rom[253][36] = -8'd41;
        rom[253][37] = -8'd1;
        rom[253][38] = 8'd10;
        rom[253][39] = -8'd7;
        rom[253][40] = 8'd19;
        rom[253][41] = -8'd3;
        rom[253][42] = -8'd1;
        rom[253][43] = -8'd1;
        rom[253][44] = 8'd12;
        rom[253][45] = -8'd3;
        rom[253][46] = 8'd7;
        rom[253][47] = 8'd30;
        rom[253][48] = -8'd21;
        rom[253][49] = 8'd5;
        rom[253][50] = -8'd10;
        rom[253][51] = -8'd10;
        rom[253][52] = 8'd42;
        rom[253][53] = 8'd19;
        rom[253][54] = 8'd18;
        rom[253][55] = -8'd22;
        rom[253][56] = 8'd15;
        rom[253][57] = 8'd1;
        rom[253][58] = 8'd5;
        rom[253][59] = 8'd13;
        rom[253][60] = -8'd2;
        rom[253][61] = -8'd15;
        rom[253][62] = -8'd25;
        rom[253][63] = -8'd20;
        rom[254][0] = 8'd8;
        rom[254][1] = -8'd11;
        rom[254][2] = -8'd24;
        rom[254][3] = 8'd28;
        rom[254][4] = -8'd19;
        rom[254][5] = 8'd16;
        rom[254][6] = -8'd11;
        rom[254][7] = 8'd1;
        rom[254][8] = 8'd0;
        rom[254][9] = -8'd7;
        rom[254][10] = 8'd21;
        rom[254][11] = 8'd28;
        rom[254][12] = -8'd5;
        rom[254][13] = -8'd22;
        rom[254][14] = -8'd42;
        rom[254][15] = 8'd39;
        rom[254][16] = 8'd27;
        rom[254][17] = 8'd40;
        rom[254][18] = 8'd32;
        rom[254][19] = -8'd38;
        rom[254][20] = -8'd14;
        rom[254][21] = -8'd2;
        rom[254][22] = -8'd55;
        rom[254][23] = -8'd29;
        rom[254][24] = -8'd31;
        rom[254][25] = 8'd40;
        rom[254][26] = -8'd22;
        rom[254][27] = 8'd0;
        rom[254][28] = -8'd13;
        rom[254][29] = -8'd24;
        rom[254][30] = -8'd85;
        rom[254][31] = 8'd6;
        rom[254][32] = -8'd4;
        rom[254][33] = -8'd33;
        rom[254][34] = 8'd13;
        rom[254][35] = -8'd5;
        rom[254][36] = 8'd12;
        rom[254][37] = -8'd2;
        rom[254][38] = -8'd46;
        rom[254][39] = -8'd35;
        rom[254][40] = -8'd11;
        rom[254][41] = -8'd30;
        rom[254][42] = -8'd35;
        rom[254][43] = -8'd64;
        rom[254][44] = 8'd24;
        rom[254][45] = -8'd6;
        rom[254][46] = 8'd1;
        rom[254][47] = 8'd16;
        rom[254][48] = -8'd3;
        rom[254][49] = -8'd50;
        rom[254][50] = -8'd15;
        rom[254][51] = 8'd37;
        rom[254][52] = -8'd47;
        rom[254][53] = 8'd18;
        rom[254][54] = 8'd27;
        rom[254][55] = -8'd33;
        rom[254][56] = -8'd29;
        rom[254][57] = -8'd18;
        rom[254][58] = -8'd9;
        rom[254][59] = -8'd10;
        rom[254][60] = 8'd18;
        rom[254][61] = -8'd9;
        rom[254][62] = 8'd23;
        rom[254][63] = 8'd12;
        rom[255][0] = -8'd67;
        rom[255][1] = 8'd16;
        rom[255][2] = -8'd2;
        rom[255][3] = -8'd11;
        rom[255][4] = 8'd15;
        rom[255][5] = 8'd5;
        rom[255][6] = 8'd23;
        rom[255][7] = 8'd17;
        rom[255][8] = -8'd38;
        rom[255][9] = -8'd18;
        rom[255][10] = 8'd3;
        rom[255][11] = 8'd4;
        rom[255][12] = -8'd16;
        rom[255][13] = -8'd6;
        rom[255][14] = -8'd16;
        rom[255][15] = 8'd33;
        rom[255][16] = -8'd3;
        rom[255][17] = -8'd37;
        rom[255][18] = -8'd21;
        rom[255][19] = -8'd33;
        rom[255][20] = -8'd2;
        rom[255][21] = -8'd4;
        rom[255][22] = -8'd3;
        rom[255][23] = 8'd17;
        rom[255][24] = 8'd38;
        rom[255][25] = -8'd14;
        rom[255][26] = 8'd11;
        rom[255][27] = -8'd43;
        rom[255][28] = -8'd9;
        rom[255][29] = -8'd60;
        rom[255][30] = -8'd42;
        rom[255][31] = -8'd11;
        rom[255][32] = 8'd16;
        rom[255][33] = -8'd6;
        rom[255][34] = -8'd59;
        rom[255][35] = 8'd23;
        rom[255][36] = -8'd20;
        rom[255][37] = 8'd46;
        rom[255][38] = -8'd34;
        rom[255][39] = 8'd16;
        rom[255][40] = -8'd33;
        rom[255][41] = 8'd18;
        rom[255][42] = 8'd16;
        rom[255][43] = -8'd26;
        rom[255][44] = 8'd19;
        rom[255][45] = 8'd21;
        rom[255][46] = 8'd1;
        rom[255][47] = 8'd20;
        rom[255][48] = -8'd46;
        rom[255][49] = 8'd46;
        rom[255][50] = -8'd17;
        rom[255][51] = -8'd6;
        rom[255][52] = 8'd10;
        rom[255][53] = 8'd9;
        rom[255][54] = -8'd17;
        rom[255][55] = -8'd24;
        rom[255][56] = 8'd0;
        rom[255][57] = -8'd30;
        rom[255][58] = 8'd0;
        rom[255][59] = -8'd20;
        rom[255][60] = 8'd6;
        rom[255][61] = 8'd3;
        rom[255][62] = -8'd17;
        rom[255][63] = -8'd8;
        rom[256][0] = -8'd16;
        rom[256][1] = 8'd14;
        rom[256][2] = -8'd24;
        rom[256][3] = -8'd16;
        rom[256][4] = -8'd33;
        rom[256][5] = -8'd16;
        rom[256][6] = -8'd16;
        rom[256][7] = -8'd7;
        rom[256][8] = -8'd25;
        rom[256][9] = 8'd17;
        rom[256][10] = 8'd3;
        rom[256][11] = 8'd20;
        rom[256][12] = 8'd9;
        rom[256][13] = -8'd10;
        rom[256][14] = 8'd16;
        rom[256][15] = 8'd11;
        rom[256][16] = 8'd4;
        rom[256][17] = -8'd1;
        rom[256][18] = 8'd17;
        rom[256][19] = -8'd5;
        rom[256][20] = 8'd5;
        rom[256][21] = -8'd49;
        rom[256][22] = -8'd40;
        rom[256][23] = -8'd26;
        rom[256][24] = 8'd9;
        rom[256][25] = -8'd14;
        rom[256][26] = -8'd20;
        rom[256][27] = 8'd0;
        rom[256][28] = -8'd14;
        rom[256][29] = -8'd11;
        rom[256][30] = 8'd35;
        rom[256][31] = -8'd22;
        rom[256][32] = -8'd9;
        rom[256][33] = -8'd24;
        rom[256][34] = -8'd15;
        rom[256][35] = -8'd24;
        rom[256][36] = -8'd39;
        rom[256][37] = 8'd24;
        rom[256][38] = -8'd8;
        rom[256][39] = 8'd2;
        rom[256][40] = -8'd3;
        rom[256][41] = -8'd24;
        rom[256][42] = 8'd2;
        rom[256][43] = 8'd8;
        rom[256][44] = -8'd26;
        rom[256][45] = 8'd27;
        rom[256][46] = 8'd7;
        rom[256][47] = -8'd8;
        rom[256][48] = 8'd8;
        rom[256][49] = 8'd29;
        rom[256][50] = -8'd4;
        rom[256][51] = -8'd52;
        rom[256][52] = 8'd5;
        rom[256][53] = -8'd22;
        rom[256][54] = -8'd11;
        rom[256][55] = 8'd31;
        rom[256][56] = -8'd30;
        rom[256][57] = -8'd4;
        rom[256][58] = 8'd21;
        rom[256][59] = 8'd28;
        rom[256][60] = -8'd21;
        rom[256][61] = 8'd6;
        rom[256][62] = -8'd11;
        rom[256][63] = -8'd9;
        rom[257][0] = -8'd56;
        rom[257][1] = -8'd57;
        rom[257][2] = -8'd23;
        rom[257][3] = 8'd13;
        rom[257][4] = -8'd27;
        rom[257][5] = -8'd41;
        rom[257][6] = -8'd20;
        rom[257][7] = -8'd47;
        rom[257][8] = 8'd11;
        rom[257][9] = 8'd15;
        rom[257][10] = -8'd49;
        rom[257][11] = -8'd14;
        rom[257][12] = -8'd44;
        rom[257][13] = -8'd60;
        rom[257][14] = -8'd12;
        rom[257][15] = -8'd56;
        rom[257][16] = -8'd1;
        rom[257][17] = 8'd14;
        rom[257][18] = -8'd27;
        rom[257][19] = -8'd60;
        rom[257][20] = -8'd23;
        rom[257][21] = -8'd9;
        rom[257][22] = -8'd31;
        rom[257][23] = -8'd43;
        rom[257][24] = -8'd14;
        rom[257][25] = 8'd18;
        rom[257][26] = -8'd10;
        rom[257][27] = -8'd94;
        rom[257][28] = 8'd10;
        rom[257][29] = 8'd17;
        rom[257][30] = 8'd11;
        rom[257][31] = -8'd23;
        rom[257][32] = -8'd51;
        rom[257][33] = -8'd25;
        rom[257][34] = -8'd32;
        rom[257][35] = 8'd2;
        rom[257][36] = -8'd24;
        rom[257][37] = -8'd41;
        rom[257][38] = 8'd3;
        rom[257][39] = 8'd19;
        rom[257][40] = 8'd15;
        rom[257][41] = -8'd31;
        rom[257][42] = -8'd24;
        rom[257][43] = -8'd41;
        rom[257][44] = 8'd1;
        rom[257][45] = -8'd70;
        rom[257][46] = -8'd30;
        rom[257][47] = -8'd1;
        rom[257][48] = -8'd42;
        rom[257][49] = 8'd6;
        rom[257][50] = -8'd94;
        rom[257][51] = 8'd5;
        rom[257][52] = 8'd5;
        rom[257][53] = -8'd65;
        rom[257][54] = 8'd10;
        rom[257][55] = -8'd52;
        rom[257][56] = -8'd1;
        rom[257][57] = 8'd34;
        rom[257][58] = 8'd32;
        rom[257][59] = -8'd26;
        rom[257][60] = -8'd9;
        rom[257][61] = -8'd24;
        rom[257][62] = -8'd13;
        rom[257][63] = 8'd25;
        rom[258][0] = -8'd44;
        rom[258][1] = -8'd24;
        rom[258][2] = -8'd23;
        rom[258][3] = -8'd41;
        rom[258][4] = -8'd65;
        rom[258][5] = 8'd0;
        rom[258][6] = -8'd14;
        rom[258][7] = 8'd0;
        rom[258][8] = -8'd21;
        rom[258][9] = 8'd34;
        rom[258][10] = 8'd18;
        rom[258][11] = -8'd40;
        rom[258][12] = 8'd0;
        rom[258][13] = 8'd20;
        rom[258][14] = -8'd21;
        rom[258][15] = -8'd11;
        rom[258][16] = -8'd36;
        rom[258][17] = 8'd14;
        rom[258][18] = 8'd15;
        rom[258][19] = -8'd34;
        rom[258][20] = -8'd12;
        rom[258][21] = -8'd19;
        rom[258][22] = -8'd24;
        rom[258][23] = -8'd15;
        rom[258][24] = 8'd16;
        rom[258][25] = -8'd12;
        rom[258][26] = -8'd12;
        rom[258][27] = -8'd6;
        rom[258][28] = 8'd12;
        rom[258][29] = -8'd13;
        rom[258][30] = -8'd1;
        rom[258][31] = -8'd41;
        rom[258][32] = -8'd45;
        rom[258][33] = -8'd25;
        rom[258][34] = -8'd7;
        rom[258][35] = -8'd22;
        rom[258][36] = 8'd0;
        rom[258][37] = -8'd1;
        rom[258][38] = -8'd4;
        rom[258][39] = -8'd10;
        rom[258][40] = -8'd59;
        rom[258][41] = -8'd27;
        rom[258][42] = -8'd59;
        rom[258][43] = -8'd28;
        rom[258][44] = -8'd8;
        rom[258][45] = -8'd3;
        rom[258][46] = -8'd44;
        rom[258][47] = -8'd22;
        rom[258][48] = -8'd3;
        rom[258][49] = 8'd9;
        rom[258][50] = -8'd29;
        rom[258][51] = 8'd17;
        rom[258][52] = 8'd43;
        rom[258][53] = -8'd49;
        rom[258][54] = -8'd44;
        rom[258][55] = 8'd6;
        rom[258][56] = -8'd19;
        rom[258][57] = -8'd20;
        rom[258][58] = -8'd26;
        rom[258][59] = -8'd11;
        rom[258][60] = -8'd2;
        rom[258][61] = 8'd19;
        rom[258][62] = 8'd25;
        rom[258][63] = -8'd39;
        rom[259][0] = 8'd0;
        rom[259][1] = 8'd30;
        rom[259][2] = 8'd21;
        rom[259][3] = 8'd36;
        rom[259][4] = 8'd3;
        rom[259][5] = 8'd3;
        rom[259][6] = 8'd51;
        rom[259][7] = 8'd19;
        rom[259][8] = -8'd3;
        rom[259][9] = -8'd2;
        rom[259][10] = -8'd39;
        rom[259][11] = -8'd8;
        rom[259][12] = -8'd42;
        rom[259][13] = 8'd16;
        rom[259][14] = -8'd13;
        rom[259][15] = 8'd27;
        rom[259][16] = -8'd23;
        rom[259][17] = -8'd41;
        rom[259][18] = 8'd19;
        rom[259][19] = 8'd24;
        rom[259][20] = -8'd4;
        rom[259][21] = 8'd29;
        rom[259][22] = 8'd25;
        rom[259][23] = 8'd8;
        rom[259][24] = 8'd13;
        rom[259][25] = 8'd24;
        rom[259][26] = -8'd15;
        rom[259][27] = 8'd1;
        rom[259][28] = -8'd7;
        rom[259][29] = -8'd5;
        rom[259][30] = 8'd10;
        rom[259][31] = -8'd12;
        rom[259][32] = -8'd6;
        rom[259][33] = -8'd12;
        rom[259][34] = -8'd36;
        rom[259][35] = 8'd8;
        rom[259][36] = 8'd9;
        rom[259][37] = 8'd15;
        rom[259][38] = 8'd40;
        rom[259][39] = 8'd27;
        rom[259][40] = 8'd1;
        rom[259][41] = -8'd7;
        rom[259][42] = 8'd35;
        rom[259][43] = 8'd5;
        rom[259][44] = 8'd4;
        rom[259][45] = -8'd38;
        rom[259][46] = 8'd12;
        rom[259][47] = -8'd41;
        rom[259][48] = 8'd11;
        rom[259][49] = 8'd13;
        rom[259][50] = -8'd11;
        rom[259][51] = -8'd8;
        rom[259][52] = 8'd18;
        rom[259][53] = -8'd6;
        rom[259][54] = -8'd30;
        rom[259][55] = -8'd18;
        rom[259][56] = 8'd20;
        rom[259][57] = -8'd60;
        rom[259][58] = -8'd11;
        rom[259][59] = -8'd2;
        rom[259][60] = 8'd18;
        rom[259][61] = -8'd5;
        rom[259][62] = 8'd4;
        rom[259][63] = 8'd29;
        rom[260][0] = -8'd14;
        rom[260][1] = -8'd22;
        rom[260][2] = -8'd8;
        rom[260][3] = -8'd4;
        rom[260][4] = -8'd15;
        rom[260][5] = -8'd9;
        rom[260][6] = -8'd4;
        rom[260][7] = -8'd16;
        rom[260][8] = 8'd13;
        rom[260][9] = -8'd4;
        rom[260][10] = -8'd31;
        rom[260][11] = -8'd24;
        rom[260][12] = -8'd61;
        rom[260][13] = -8'd22;
        rom[260][14] = 8'd4;
        rom[260][15] = 8'd27;
        rom[260][16] = 8'd22;
        rom[260][17] = 8'd0;
        rom[260][18] = 8'd33;
        rom[260][19] = 8'd10;
        rom[260][20] = -8'd2;
        rom[260][21] = -8'd40;
        rom[260][22] = 8'd12;
        rom[260][23] = 8'd26;
        rom[260][24] = -8'd40;
        rom[260][25] = -8'd7;
        rom[260][26] = -8'd17;
        rom[260][27] = -8'd5;
        rom[260][28] = -8'd32;
        rom[260][29] = -8'd3;
        rom[260][30] = -8'd41;
        rom[260][31] = -8'd16;
        rom[260][32] = 8'd3;
        rom[260][33] = 8'd36;
        rom[260][34] = -8'd30;
        rom[260][35] = -8'd7;
        rom[260][36] = -8'd23;
        rom[260][37] = 8'd2;
        rom[260][38] = -8'd51;
        rom[260][39] = -8'd3;
        rom[260][40] = -8'd21;
        rom[260][41] = -8'd25;
        rom[260][42] = 8'd8;
        rom[260][43] = -8'd32;
        rom[260][44] = -8'd20;
        rom[260][45] = -8'd42;
        rom[260][46] = -8'd49;
        rom[260][47] = -8'd5;
        rom[260][48] = 8'd3;
        rom[260][49] = -8'd10;
        rom[260][50] = -8'd18;
        rom[260][51] = -8'd24;
        rom[260][52] = -8'd44;
        rom[260][53] = -8'd17;
        rom[260][54] = -8'd8;
        rom[260][55] = 8'd5;
        rom[260][56] = -8'd7;
        rom[260][57] = -8'd15;
        rom[260][58] = 8'd25;
        rom[260][59] = -8'd8;
        rom[260][60] = 8'd10;
        rom[260][61] = 8'd28;
        rom[260][62] = 8'd5;
        rom[260][63] = -8'd50;
        rom[261][0] = -8'd1;
        rom[261][1] = 8'd2;
        rom[261][2] = -8'd4;
        rom[261][3] = -8'd5;
        rom[261][4] = -8'd7;
        rom[261][5] = 8'd14;
        rom[261][6] = -8'd5;
        rom[261][7] = 8'd11;
        rom[261][8] = -8'd5;
        rom[261][9] = 8'd3;
        rom[261][10] = -8'd6;
        rom[261][11] = 8'd2;
        rom[261][12] = -8'd3;
        rom[261][13] = 8'd3;
        rom[261][14] = 8'd7;
        rom[261][15] = 8'd1;
        rom[261][16] = 8'd2;
        rom[261][17] = -8'd7;
        rom[261][18] = -8'd5;
        rom[261][19] = 8'd0;
        rom[261][20] = 8'd8;
        rom[261][21] = 8'd7;
        rom[261][22] = 8'd12;
        rom[261][23] = 8'd10;
        rom[261][24] = 8'd11;
        rom[261][25] = -8'd12;
        rom[261][26] = 8'd0;
        rom[261][27] = -8'd4;
        rom[261][28] = -8'd4;
        rom[261][29] = -8'd6;
        rom[261][30] = -8'd15;
        rom[261][31] = -8'd8;
        rom[261][32] = -8'd9;
        rom[261][33] = 8'd1;
        rom[261][34] = 8'd4;
        rom[261][35] = -8'd8;
        rom[261][36] = 8'd5;
        rom[261][37] = 8'd5;
        rom[261][38] = -8'd2;
        rom[261][39] = 8'd3;
        rom[261][40] = 8'd5;
        rom[261][41] = -8'd7;
        rom[261][42] = -8'd3;
        rom[261][43] = 8'd1;
        rom[261][44] = -8'd4;
        rom[261][45] = 8'd4;
        rom[261][46] = -8'd3;
        rom[261][47] = 8'd10;
        rom[261][48] = -8'd6;
        rom[261][49] = -8'd5;
        rom[261][50] = -8'd2;
        rom[261][51] = 8'd4;
        rom[261][52] = 8'd4;
        rom[261][53] = 8'd10;
        rom[261][54] = 8'd9;
        rom[261][55] = -8'd7;
        rom[261][56] = 8'd12;
        rom[261][57] = -8'd6;
        rom[261][58] = 8'd6;
        rom[261][59] = -8'd5;
        rom[261][60] = 8'd1;
        rom[261][61] = 8'd6;
        rom[261][62] = 8'd1;
        rom[261][63] = -8'd7;
        rom[262][0] = 8'd12;
        rom[262][1] = -8'd42;
        rom[262][2] = 8'd31;
        rom[262][3] = 8'd24;
        rom[262][4] = -8'd36;
        rom[262][5] = 8'd4;
        rom[262][6] = -8'd24;
        rom[262][7] = -8'd11;
        rom[262][8] = 8'd9;
        rom[262][9] = 8'd33;
        rom[262][10] = -8'd25;
        rom[262][11] = 8'd35;
        rom[262][12] = -8'd14;
        rom[262][13] = 8'd8;
        rom[262][14] = 8'd7;
        rom[262][15] = -8'd14;
        rom[262][16] = -8'd44;
        rom[262][17] = 8'd3;
        rom[262][18] = 8'd1;
        rom[262][19] = -8'd3;
        rom[262][20] = 8'd4;
        rom[262][21] = -8'd58;
        rom[262][22] = 8'd5;
        rom[262][23] = 8'd17;
        rom[262][24] = 8'd1;
        rom[262][25] = -8'd19;
        rom[262][26] = 8'd3;
        rom[262][27] = -8'd1;
        rom[262][28] = 8'd33;
        rom[262][29] = 8'd3;
        rom[262][30] = -8'd5;
        rom[262][31] = 8'd14;
        rom[262][32] = -8'd39;
        rom[262][33] = 8'd22;
        rom[262][34] = 8'd0;
        rom[262][35] = -8'd37;
        rom[262][36] = -8'd2;
        rom[262][37] = -8'd6;
        rom[262][38] = 8'd10;
        rom[262][39] = -8'd9;
        rom[262][40] = -8'd42;
        rom[262][41] = -8'd21;
        rom[262][42] = 8'd17;
        rom[262][43] = -8'd21;
        rom[262][44] = 8'd0;
        rom[262][45] = -8'd9;
        rom[262][46] = -8'd39;
        rom[262][47] = -8'd47;
        rom[262][48] = 8'd53;
        rom[262][49] = -8'd9;
        rom[262][50] = 8'd5;
        rom[262][51] = -8'd14;
        rom[262][52] = -8'd9;
        rom[262][53] = 8'd16;
        rom[262][54] = 8'd23;
        rom[262][55] = -8'd23;
        rom[262][56] = -8'd34;
        rom[262][57] = 8'd33;
        rom[262][58] = -8'd9;
        rom[262][59] = -8'd37;
        rom[262][60] = -8'd6;
        rom[262][61] = -8'd9;
        rom[262][62] = -8'd5;
        rom[262][63] = -8'd7;
        rom[263][0] = 8'd8;
        rom[263][1] = -8'd24;
        rom[263][2] = -8'd77;
        rom[263][3] = 8'd3;
        rom[263][4] = -8'd46;
        rom[263][5] = -8'd29;
        rom[263][6] = 8'd3;
        rom[263][7] = 8'd9;
        rom[263][8] = -8'd14;
        rom[263][9] = -8'd21;
        rom[263][10] = -8'd5;
        rom[263][11] = -8'd5;
        rom[263][12] = -8'd10;
        rom[263][13] = 8'd2;
        rom[263][14] = -8'd37;
        rom[263][15] = 8'd15;
        rom[263][16] = -8'd12;
        rom[263][17] = 8'd30;
        rom[263][18] = -8'd28;
        rom[263][19] = 8'd10;
        rom[263][20] = -8'd8;
        rom[263][21] = 8'd25;
        rom[263][22] = 8'd3;
        rom[263][23] = 8'd29;
        rom[263][24] = -8'd14;
        rom[263][25] = -8'd3;
        rom[263][26] = 8'd1;
        rom[263][27] = -8'd5;
        rom[263][28] = 8'd36;
        rom[263][29] = 8'd13;
        rom[263][30] = -8'd49;
        rom[263][31] = -8'd4;
        rom[263][32] = -8'd16;
        rom[263][33] = 8'd31;
        rom[263][34] = 8'd10;
        rom[263][35] = -8'd76;
        rom[263][36] = -8'd43;
        rom[263][37] = -8'd26;
        rom[263][38] = 8'd14;
        rom[263][39] = 8'd4;
        rom[263][40] = 8'd11;
        rom[263][41] = -8'd20;
        rom[263][42] = 8'd14;
        rom[263][43] = 8'd25;
        rom[263][44] = 8'd14;
        rom[263][45] = 8'd35;
        rom[263][46] = 8'd27;
        rom[263][47] = 8'd48;
        rom[263][48] = -8'd35;
        rom[263][49] = 8'd24;
        rom[263][50] = -8'd31;
        rom[263][51] = 8'd1;
        rom[263][52] = -8'd28;
        rom[263][53] = -8'd37;
        rom[263][54] = -8'd75;
        rom[263][55] = -8'd3;
        rom[263][56] = 8'd13;
        rom[263][57] = 8'd1;
        rom[263][58] = -8'd10;
        rom[263][59] = -8'd21;
        rom[263][60] = -8'd6;
        rom[263][61] = -8'd28;
        rom[263][62] = 8'd17;
        rom[263][63] = 8'd19;
        rom[264][0] = 8'd10;
        rom[264][1] = 8'd1;
        rom[264][2] = 8'd9;
        rom[264][3] = 8'd7;
        rom[264][4] = 8'd8;
        rom[264][5] = -8'd16;
        rom[264][6] = -8'd21;
        rom[264][7] = -8'd27;
        rom[264][8] = -8'd2;
        rom[264][9] = -8'd12;
        rom[264][10] = 8'd9;
        rom[264][11] = -8'd66;
        rom[264][12] = -8'd7;
        rom[264][13] = -8'd6;
        rom[264][14] = -8'd22;
        rom[264][15] = 8'd2;
        rom[264][16] = 8'd6;
        rom[264][17] = -8'd18;
        rom[264][18] = -8'd25;
        rom[264][19] = 8'd13;
        rom[264][20] = -8'd16;
        rom[264][21] = 8'd13;
        rom[264][22] = -8'd21;
        rom[264][23] = 8'd8;
        rom[264][24] = -8'd40;
        rom[264][25] = 8'd9;
        rom[264][26] = -8'd12;
        rom[264][27] = -8'd15;
        rom[264][28] = 8'd6;
        rom[264][29] = 8'd12;
        rom[264][30] = -8'd64;
        rom[264][31] = 8'd8;
        rom[264][32] = 8'd13;
        rom[264][33] = 8'd18;
        rom[264][34] = -8'd15;
        rom[264][35] = -8'd21;
        rom[264][36] = -8'd16;
        rom[264][37] = 8'd0;
        rom[264][38] = -8'd35;
        rom[264][39] = -8'd19;
        rom[264][40] = -8'd14;
        rom[264][41] = -8'd6;
        rom[264][42] = 8'd15;
        rom[264][43] = 8'd7;
        rom[264][44] = 8'd30;
        rom[264][45] = -8'd22;
        rom[264][46] = 8'd6;
        rom[264][47] = 8'd1;
        rom[264][48] = -8'd3;
        rom[264][49] = -8'd8;
        rom[264][50] = -8'd14;
        rom[264][51] = -8'd26;
        rom[264][52] = -8'd2;
        rom[264][53] = -8'd39;
        rom[264][54] = -8'd7;
        rom[264][55] = -8'd4;
        rom[264][56] = 8'd8;
        rom[264][57] = -8'd31;
        rom[264][58] = -8'd6;
        rom[264][59] = -8'd26;
        rom[264][60] = -8'd8;
        rom[264][61] = -8'd37;
        rom[264][62] = -8'd5;
        rom[264][63] = -8'd39;
        rom[265][0] = -8'd45;
        rom[265][1] = -8'd17;
        rom[265][2] = 8'd14;
        rom[265][3] = -8'd9;
        rom[265][4] = 8'd12;
        rom[265][5] = 8'd18;
        rom[265][6] = -8'd36;
        rom[265][7] = 8'd26;
        rom[265][8] = -8'd33;
        rom[265][9] = -8'd6;
        rom[265][10] = -8'd12;
        rom[265][11] = -8'd11;
        rom[265][12] = 8'd5;
        rom[265][13] = 8'd9;
        rom[265][14] = 8'd32;
        rom[265][15] = -8'd39;
        rom[265][16] = -8'd16;
        rom[265][17] = 8'd21;
        rom[265][18] = 8'd15;
        rom[265][19] = -8'd21;
        rom[265][20] = -8'd4;
        rom[265][21] = -8'd17;
        rom[265][22] = 8'd27;
        rom[265][23] = -8'd9;
        rom[265][24] = -8'd10;
        rom[265][25] = -8'd9;
        rom[265][26] = 8'd4;
        rom[265][27] = -8'd11;
        rom[265][28] = -8'd21;
        rom[265][29] = -8'd12;
        rom[265][30] = -8'd26;
        rom[265][31] = 8'd22;
        rom[265][32] = 8'd2;
        rom[265][33] = -8'd25;
        rom[265][34] = 8'd25;
        rom[265][35] = 8'd10;
        rom[265][36] = -8'd57;
        rom[265][37] = 8'd18;
        rom[265][38] = 8'd28;
        rom[265][39] = -8'd38;
        rom[265][40] = -8'd18;
        rom[265][41] = -8'd43;
        rom[265][42] = 8'd64;
        rom[265][43] = 8'd8;
        rom[265][44] = 8'd18;
        rom[265][45] = -8'd5;
        rom[265][46] = -8'd6;
        rom[265][47] = 8'd16;
        rom[265][48] = 8'd24;
        rom[265][49] = -8'd25;
        rom[265][50] = 8'd5;
        rom[265][51] = -8'd14;
        rom[265][52] = 8'd20;
        rom[265][53] = 8'd35;
        rom[265][54] = -8'd29;
        rom[265][55] = 8'd22;
        rom[265][56] = 8'd2;
        rom[265][57] = -8'd9;
        rom[265][58] = 8'd15;
        rom[265][59] = 8'd35;
        rom[265][60] = 8'd17;
        rom[265][61] = 8'd27;
        rom[265][62] = 8'd18;
        rom[265][63] = -8'd3;
        rom[266][0] = 8'd4;
        rom[266][1] = 8'd0;
        rom[266][2] = 8'd11;
        rom[266][3] = -8'd13;
        rom[266][4] = -8'd11;
        rom[266][5] = -8'd8;
        rom[266][6] = 8'd5;
        rom[266][7] = -8'd5;
        rom[266][8] = 8'd4;
        rom[266][9] = -8'd18;
        rom[266][10] = 8'd33;
        rom[266][11] = 8'd8;
        rom[266][12] = 8'd30;
        rom[266][13] = 8'd36;
        rom[266][14] = -8'd14;
        rom[266][15] = 8'd15;
        rom[266][16] = -8'd25;
        rom[266][17] = -8'd15;
        rom[266][18] = -8'd28;
        rom[266][19] = 8'd11;
        rom[266][20] = -8'd5;
        rom[266][21] = 8'd14;
        rom[266][22] = -8'd7;
        rom[266][23] = -8'd47;
        rom[266][24] = 8'd25;
        rom[266][25] = 8'd20;
        rom[266][26] = -8'd22;
        rom[266][27] = 8'd56;
        rom[266][28] = -8'd20;
        rom[266][29] = 8'd0;
        rom[266][30] = 8'd16;
        rom[266][31] = 8'd22;
        rom[266][32] = 8'd9;
        rom[266][33] = -8'd19;
        rom[266][34] = -8'd4;
        rom[266][35] = -8'd12;
        rom[266][36] = 8'd3;
        rom[266][37] = 8'd12;
        rom[266][38] = 8'd30;
        rom[266][39] = 8'd3;
        rom[266][40] = 8'd11;
        rom[266][41] = 8'd1;
        rom[266][42] = -8'd7;
        rom[266][43] = -8'd14;
        rom[266][44] = 8'd22;
        rom[266][45] = 8'd24;
        rom[266][46] = -8'd4;
        rom[266][47] = 8'd6;
        rom[266][48] = 8'd7;
        rom[266][49] = 8'd22;
        rom[266][50] = -8'd10;
        rom[266][51] = 8'd5;
        rom[266][52] = -8'd14;
        rom[266][53] = -8'd1;
        rom[266][54] = -8'd18;
        rom[266][55] = -8'd21;
        rom[266][56] = -8'd38;
        rom[266][57] = -8'd3;
        rom[266][58] = 8'd24;
        rom[266][59] = -8'd8;
        rom[266][60] = 8'd5;
        rom[266][61] = -8'd31;
        rom[266][62] = -8'd37;
        rom[266][63] = -8'd11;
        rom[267][0] = -8'd45;
        rom[267][1] = 8'd16;
        rom[267][2] = 8'd16;
        rom[267][3] = -8'd35;
        rom[267][4] = 8'd14;
        rom[267][5] = 8'd8;
        rom[267][6] = 8'd13;
        rom[267][7] = -8'd6;
        rom[267][8] = -8'd7;
        rom[267][9] = 8'd4;
        rom[267][10] = -8'd10;
        rom[267][11] = -8'd14;
        rom[267][12] = 8'd2;
        rom[267][13] = 8'd44;
        rom[267][14] = -8'd6;
        rom[267][15] = -8'd8;
        rom[267][16] = 8'd13;
        rom[267][17] = -8'd7;
        rom[267][18] = -8'd6;
        rom[267][19] = 8'd9;
        rom[267][20] = 8'd2;
        rom[267][21] = 8'd21;
        rom[267][22] = 8'd18;
        rom[267][23] = 8'd12;
        rom[267][24] = 8'd14;
        rom[267][25] = -8'd41;
        rom[267][26] = 8'd15;
        rom[267][27] = 8'd7;
        rom[267][28] = 8'd44;
        rom[267][29] = 8'd43;
        rom[267][30] = 8'd33;
        rom[267][31] = -8'd42;
        rom[267][32] = -8'd37;
        rom[267][33] = 8'd12;
        rom[267][34] = 8'd15;
        rom[267][35] = 8'd6;
        rom[267][36] = -8'd18;
        rom[267][37] = -8'd41;
        rom[267][38] = -8'd17;
        rom[267][39] = -8'd8;
        rom[267][40] = -8'd18;
        rom[267][41] = -8'd4;
        rom[267][42] = 8'd9;
        rom[267][43] = -8'd13;
        rom[267][44] = -8'd45;
        rom[267][45] = -8'd2;
        rom[267][46] = 8'd27;
        rom[267][47] = 8'd19;
        rom[267][48] = 8'd7;
        rom[267][49] = -8'd42;
        rom[267][50] = -8'd32;
        rom[267][51] = 8'd49;
        rom[267][52] = -8'd45;
        rom[267][53] = -8'd57;
        rom[267][54] = -8'd2;
        rom[267][55] = -8'd43;
        rom[267][56] = -8'd16;
        rom[267][57] = -8'd23;
        rom[267][58] = 8'd9;
        rom[267][59] = 8'd13;
        rom[267][60] = -8'd58;
        rom[267][61] = -8'd7;
        rom[267][62] = 8'd5;
        rom[267][63] = -8'd3;
        rom[268][0] = -8'd71;
        rom[268][1] = -8'd42;
        rom[268][2] = 8'd46;
        rom[268][3] = 8'd17;
        rom[268][4] = 8'd6;
        rom[268][5] = -8'd55;
        rom[268][6] = 8'd6;
        rom[268][7] = -8'd67;
        rom[268][8] = -8'd3;
        rom[268][9] = 8'd22;
        rom[268][10] = 8'd24;
        rom[268][11] = -8'd10;
        rom[268][12] = -8'd48;
        rom[268][13] = 8'd3;
        rom[268][14] = 8'd11;
        rom[268][15] = 8'd35;
        rom[268][16] = 8'd9;
        rom[268][17] = -8'd36;
        rom[268][18] = 8'd0;
        rom[268][19] = -8'd94;
        rom[268][20] = -8'd1;
        rom[268][21] = 8'd3;
        rom[268][22] = -8'd18;
        rom[268][23] = -8'd33;
        rom[268][24] = -8'd7;
        rom[268][25] = 8'd13;
        rom[268][26] = -8'd16;
        rom[268][27] = -8'd7;
        rom[268][28] = 8'd2;
        rom[268][29] = -8'd8;
        rom[268][30] = -8'd14;
        rom[268][31] = 8'd5;
        rom[268][32] = 8'd17;
        rom[268][33] = 8'd11;
        rom[268][34] = 8'd6;
        rom[268][35] = -8'd19;
        rom[268][36] = -8'd21;
        rom[268][37] = -8'd30;
        rom[268][38] = 8'd18;
        rom[268][39] = -8'd4;
        rom[268][40] = -8'd43;
        rom[268][41] = -8'd4;
        rom[268][42] = -8'd23;
        rom[268][43] = 8'd4;
        rom[268][44] = -8'd9;
        rom[268][45] = -8'd61;
        rom[268][46] = -8'd13;
        rom[268][47] = 8'd54;
        rom[268][48] = -8'd3;
        rom[268][49] = 8'd24;
        rom[268][50] = 8'd15;
        rom[268][51] = -8'd1;
        rom[268][52] = -8'd49;
        rom[268][53] = -8'd6;
        rom[268][54] = 8'd19;
        rom[268][55] = 8'd11;
        rom[268][56] = -8'd20;
        rom[268][57] = 8'd38;
        rom[268][58] = -8'd34;
        rom[268][59] = -8'd1;
        rom[268][60] = 8'd4;
        rom[268][61] = -8'd1;
        rom[268][62] = 8'd5;
        rom[268][63] = 8'd24;
        rom[269][0] = 8'd39;
        rom[269][1] = -8'd8;
        rom[269][2] = 8'd24;
        rom[269][3] = -8'd35;
        rom[269][4] = 8'd22;
        rom[269][5] = 8'd52;
        rom[269][6] = -8'd21;
        rom[269][7] = 8'd20;
        rom[269][8] = -8'd13;
        rom[269][9] = 8'd8;
        rom[269][10] = -8'd6;
        rom[269][11] = -8'd19;
        rom[269][12] = 8'd1;
        rom[269][13] = 8'd18;
        rom[269][14] = 8'd20;
        rom[269][15] = 8'd12;
        rom[269][16] = 8'd0;
        rom[269][17] = -8'd40;
        rom[269][18] = -8'd3;
        rom[269][19] = 8'd11;
        rom[269][20] = 8'd4;
        rom[269][21] = -8'd9;
        rom[269][22] = -8'd24;
        rom[269][23] = 8'd15;
        rom[269][24] = -8'd16;
        rom[269][25] = -8'd47;
        rom[269][26] = -8'd5;
        rom[269][27] = 8'd7;
        rom[269][28] = -8'd11;
        rom[269][29] = 8'd45;
        rom[269][30] = 8'd18;
        rom[269][31] = -8'd7;
        rom[269][32] = -8'd1;
        rom[269][33] = 8'd8;
        rom[269][34] = -8'd49;
        rom[269][35] = -8'd20;
        rom[269][36] = -8'd7;
        rom[269][37] = -8'd22;
        rom[269][38] = -8'd3;
        rom[269][39] = 8'd4;
        rom[269][40] = -8'd20;
        rom[269][41] = -8'd1;
        rom[269][42] = -8'd26;
        rom[269][43] = 8'd0;
        rom[269][44] = 8'd10;
        rom[269][45] = -8'd19;
        rom[269][46] = -8'd19;
        rom[269][47] = -8'd50;
        rom[269][48] = 8'd5;
        rom[269][49] = -8'd34;
        rom[269][50] = 8'd16;
        rom[269][51] = -8'd43;
        rom[269][52] = 8'd9;
        rom[269][53] = 8'd32;
        rom[269][54] = 8'd6;
        rom[269][55] = 8'd12;
        rom[269][56] = 8'd8;
        rom[269][57] = 8'd0;
        rom[269][58] = 8'd20;
        rom[269][59] = 8'd12;
        rom[269][60] = -8'd19;
        rom[269][61] = -8'd1;
        rom[269][62] = 8'd14;
        rom[269][63] = 8'd9;
        rom[270][0] = 8'd14;
        rom[270][1] = 8'd6;
        rom[270][2] = 8'd30;
        rom[270][3] = -8'd27;
        rom[270][4] = 8'd15;
        rom[270][5] = -8'd22;
        rom[270][6] = 8'd8;
        rom[270][7] = -8'd72;
        rom[270][8] = -8'd13;
        rom[270][9] = -8'd49;
        rom[270][10] = 8'd16;
        rom[270][11] = -8'd30;
        rom[270][12] = -8'd3;
        rom[270][13] = 8'd13;
        rom[270][14] = -8'd14;
        rom[270][15] = -8'd14;
        rom[270][16] = -8'd6;
        rom[270][17] = -8'd36;
        rom[270][18] = -8'd34;
        rom[270][19] = -8'd20;
        rom[270][20] = -8'd8;
        rom[270][21] = 8'd10;
        rom[270][22] = -8'd2;
        rom[270][23] = 8'd16;
        rom[270][24] = -8'd13;
        rom[270][25] = -8'd21;
        rom[270][26] = 8'd2;
        rom[270][27] = 8'd25;
        rom[270][28] = -8'd60;
        rom[270][29] = -8'd22;
        rom[270][30] = -8'd16;
        rom[270][31] = -8'd7;
        rom[270][32] = -8'd13;
        rom[270][33] = 8'd36;
        rom[270][34] = 8'd17;
        rom[270][35] = 8'd9;
        rom[270][36] = 8'd19;
        rom[270][37] = 8'd14;
        rom[270][38] = -8'd42;
        rom[270][39] = 8'd29;
        rom[270][40] = -8'd2;
        rom[270][41] = -8'd22;
        rom[270][42] = 8'd0;
        rom[270][43] = 8'd6;
        rom[270][44] = -8'd11;
        rom[270][45] = -8'd44;
        rom[270][46] = 8'd29;
        rom[270][47] = -8'd45;
        rom[270][48] = 8'd3;
        rom[270][49] = -8'd22;
        rom[270][50] = -8'd9;
        rom[270][51] = 8'd19;
        rom[270][52] = -8'd13;
        rom[270][53] = -8'd9;
        rom[270][54] = 8'd23;
        rom[270][55] = -8'd32;
        rom[270][56] = -8'd5;
        rom[270][57] = 8'd1;
        rom[270][58] = 8'd17;
        rom[270][59] = 8'd4;
        rom[270][60] = -8'd18;
        rom[270][61] = 8'd5;
        rom[270][62] = 8'd32;
        rom[270][63] = -8'd18;
        rom[271][0] = 8'd1;
        rom[271][1] = -8'd49;
        rom[271][2] = -8'd4;
        rom[271][3] = 8'd3;
        rom[271][4] = 8'd8;
        rom[271][5] = 8'd7;
        rom[271][6] = 8'd0;
        rom[271][7] = -8'd36;
        rom[271][8] = 8'd7;
        rom[271][9] = 8'd10;
        rom[271][10] = -8'd22;
        rom[271][11] = -8'd6;
        rom[271][12] = 8'd32;
        rom[271][13] = -8'd12;
        rom[271][14] = 8'd7;
        rom[271][15] = -8'd15;
        rom[271][16] = -8'd19;
        rom[271][17] = 8'd28;
        rom[271][18] = 8'd12;
        rom[271][19] = -8'd15;
        rom[271][20] = 8'd1;
        rom[271][21] = -8'd23;
        rom[271][22] = -8'd5;
        rom[271][23] = -8'd3;
        rom[271][24] = -8'd66;
        rom[271][25] = -8'd2;
        rom[271][26] = -8'd9;
        rom[271][27] = 8'd5;
        rom[271][28] = 8'd9;
        rom[271][29] = -8'd16;
        rom[271][30] = -8'd20;
        rom[271][31] = -8'd34;
        rom[271][32] = -8'd31;
        rom[271][33] = -8'd1;
        rom[271][34] = 8'd20;
        rom[271][35] = 8'd23;
        rom[271][36] = 8'd4;
        rom[271][37] = 8'd3;
        rom[271][38] = -8'd16;
        rom[271][39] = 8'd9;
        rom[271][40] = -8'd19;
        rom[271][41] = -8'd2;
        rom[271][42] = 8'd6;
        rom[271][43] = -8'd11;
        rom[271][44] = 8'd11;
        rom[271][45] = -8'd18;
        rom[271][46] = 8'd12;
        rom[271][47] = -8'd4;
        rom[271][48] = 8'd31;
        rom[271][49] = -8'd22;
        rom[271][50] = -8'd7;
        rom[271][51] = -8'd28;
        rom[271][52] = 8'd0;
        rom[271][53] = 8'd18;
        rom[271][54] = 8'd10;
        rom[271][55] = -8'd49;
        rom[271][56] = 8'd14;
        rom[271][57] = -8'd24;
        rom[271][58] = -8'd33;
        rom[271][59] = 8'd17;
        rom[271][60] = 8'd15;
        rom[271][61] = -8'd33;
        rom[271][62] = -8'd32;
        rom[271][63] = 8'd12;
        rom[272][0] = 8'd7;
        rom[272][1] = -8'd4;
        rom[272][2] = 8'd7;
        rom[272][3] = 8'd3;
        rom[272][4] = 8'd5;
        rom[272][5] = -8'd7;
        rom[272][6] = 8'd5;
        rom[272][7] = 8'd2;
        rom[272][8] = 8'd10;
        rom[272][9] = 8'd3;
        rom[272][10] = -8'd3;
        rom[272][11] = -8'd6;
        rom[272][12] = 8'd4;
        rom[272][13] = 8'd0;
        rom[272][14] = -8'd7;
        rom[272][15] = -8'd7;
        rom[272][16] = -8'd6;
        rom[272][17] = -8'd1;
        rom[272][18] = 8'd0;
        rom[272][19] = 8'd6;
        rom[272][20] = 8'd0;
        rom[272][21] = 8'd2;
        rom[272][22] = -8'd2;
        rom[272][23] = -8'd8;
        rom[272][24] = 8'd3;
        rom[272][25] = 8'd6;
        rom[272][26] = -8'd4;
        rom[272][27] = -8'd3;
        rom[272][28] = 8'd10;
        rom[272][29] = -8'd6;
        rom[272][30] = -8'd5;
        rom[272][31] = 8'd7;
        rom[272][32] = -8'd6;
        rom[272][33] = -8'd5;
        rom[272][34] = -8'd4;
        rom[272][35] = 8'd5;
        rom[272][36] = -8'd4;
        rom[272][37] = -8'd5;
        rom[272][38] = 8'd7;
        rom[272][39] = -8'd3;
        rom[272][40] = -8'd5;
        rom[272][41] = -8'd8;
        rom[272][42] = -8'd1;
        rom[272][43] = 8'd7;
        rom[272][44] = 8'd2;
        rom[272][45] = 8'd0;
        rom[272][46] = -8'd4;
        rom[272][47] = 8'd6;
        rom[272][48] = 8'd8;
        rom[272][49] = 8'd0;
        rom[272][50] = -8'd1;
        rom[272][51] = -8'd11;
        rom[272][52] = 8'd4;
        rom[272][53] = 8'd5;
        rom[272][54] = 8'd7;
        rom[272][55] = -8'd3;
        rom[272][56] = -8'd4;
        rom[272][57] = 8'd1;
        rom[272][58] = 8'd2;
        rom[272][59] = -8'd2;
        rom[272][60] = -8'd3;
        rom[272][61] = 8'd8;
        rom[272][62] = -8'd7;
        rom[272][63] = 8'd1;
        rom[273][0] = -8'd58;
        rom[273][1] = 8'd58;
        rom[273][2] = -8'd15;
        rom[273][3] = -8'd6;
        rom[273][4] = -8'd10;
        rom[273][5] = -8'd25;
        rom[273][6] = 8'd3;
        rom[273][7] = 8'd15;
        rom[273][8] = 8'd40;
        rom[273][9] = 8'd23;
        rom[273][10] = -8'd53;
        rom[273][11] = 8'd12;
        rom[273][12] = 8'd21;
        rom[273][13] = -8'd15;
        rom[273][14] = -8'd6;
        rom[273][15] = -8'd29;
        rom[273][16] = 8'd11;
        rom[273][17] = 8'd23;
        rom[273][18] = 8'd10;
        rom[273][19] = -8'd23;
        rom[273][20] = -8'd6;
        rom[273][21] = -8'd23;
        rom[273][22] = -8'd6;
        rom[273][23] = -8'd28;
        rom[273][24] = 8'd7;
        rom[273][25] = 8'd2;
        rom[273][26] = -8'd33;
        rom[273][27] = -8'd50;
        rom[273][28] = -8'd23;
        rom[273][29] = -8'd1;
        rom[273][30] = 8'd14;
        rom[273][31] = 8'd12;
        rom[273][32] = 8'd18;
        rom[273][33] = 8'd6;
        rom[273][34] = -8'd14;
        rom[273][35] = -8'd21;
        rom[273][36] = 8'd9;
        rom[273][37] = 8'd23;
        rom[273][38] = -8'd3;
        rom[273][39] = 8'd24;
        rom[273][40] = -8'd14;
        rom[273][41] = 8'd25;
        rom[273][42] = 8'd22;
        rom[273][43] = 8'd8;
        rom[273][44] = 8'd31;
        rom[273][45] = 8'd9;
        rom[273][46] = -8'd27;
        rom[273][47] = 8'd3;
        rom[273][48] = -8'd45;
        rom[273][49] = 8'd12;
        rom[273][50] = 8'd24;
        rom[273][51] = 8'd3;
        rom[273][52] = 8'd7;
        rom[273][53] = 8'd20;
        rom[273][54] = -8'd5;
        rom[273][55] = -8'd4;
        rom[273][56] = 8'd0;
        rom[273][57] = -8'd19;
        rom[273][58] = -8'd14;
        rom[273][59] = 8'd11;
        rom[273][60] = 8'd7;
        rom[273][61] = 8'd34;
        rom[273][62] = -8'd48;
        rom[273][63] = -8'd40;
        rom[274][0] = 8'd35;
        rom[274][1] = 8'd0;
        rom[274][2] = 8'd19;
        rom[274][3] = -8'd17;
        rom[274][4] = -8'd23;
        rom[274][5] = 8'd11;
        rom[274][6] = 8'd7;
        rom[274][7] = 8'd13;
        rom[274][8] = 8'd15;
        rom[274][9] = 8'd4;
        rom[274][10] = -8'd12;
        rom[274][11] = -8'd5;
        rom[274][12] = 8'd11;
        rom[274][13] = 8'd12;
        rom[274][14] = 8'd13;
        rom[274][15] = -8'd29;
        rom[274][16] = -8'd55;
        rom[274][17] = -8'd29;
        rom[274][18] = -8'd1;
        rom[274][19] = -8'd4;
        rom[274][20] = -8'd7;
        rom[274][21] = -8'd46;
        rom[274][22] = 8'd23;
        rom[274][23] = 8'd7;
        rom[274][24] = 8'd16;
        rom[274][25] = -8'd49;
        rom[274][26] = -8'd25;
        rom[274][27] = 8'd31;
        rom[274][28] = -8'd16;
        rom[274][29] = -8'd17;
        rom[274][30] = -8'd3;
        rom[274][31] = 8'd4;
        rom[274][32] = -8'd11;
        rom[274][33] = 8'd40;
        rom[274][34] = 8'd1;
        rom[274][35] = -8'd12;
        rom[274][36] = 8'd6;
        rom[274][37] = -8'd21;
        rom[274][38] = -8'd50;
        rom[274][39] = 8'd23;
        rom[274][40] = 8'd1;
        rom[274][41] = 8'd21;
        rom[274][42] = 8'd18;
        rom[274][43] = -8'd39;
        rom[274][44] = -8'd4;
        rom[274][45] = 8'd21;
        rom[274][46] = -8'd26;
        rom[274][47] = -8'd76;
        rom[274][48] = -8'd11;
        rom[274][49] = 8'd8;
        rom[274][50] = 8'd10;
        rom[274][51] = -8'd13;
        rom[274][52] = -8'd13;
        rom[274][53] = -8'd11;
        rom[274][54] = 8'd16;
        rom[274][55] = 8'd9;
        rom[274][56] = 8'd14;
        rom[274][57] = -8'd39;
        rom[274][58] = -8'd67;
        rom[274][59] = -8'd31;
        rom[274][60] = -8'd10;
        rom[274][61] = -8'd42;
        rom[274][62] = 8'd23;
        rom[274][63] = 8'd17;
        rom[275][0] = -8'd33;
        rom[275][1] = -8'd39;
        rom[275][2] = -8'd53;
        rom[275][3] = -8'd65;
        rom[275][4] = 8'd11;
        rom[275][5] = -8'd2;
        rom[275][6] = -8'd43;
        rom[275][7] = -8'd5;
        rom[275][8] = -8'd36;
        rom[275][9] = -8'd4;
        rom[275][10] = -8'd27;
        rom[275][11] = -8'd44;
        rom[275][12] = 8'd3;
        rom[275][13] = 8'd7;
        rom[275][14] = 8'd14;
        rom[275][15] = -8'd22;
        rom[275][16] = -8'd3;
        rom[275][17] = -8'd18;
        rom[275][18] = -8'd35;
        rom[275][19] = -8'd38;
        rom[275][20] = 8'd0;
        rom[275][21] = -8'd59;
        rom[275][22] = -8'd39;
        rom[275][23] = -8'd35;
        rom[275][24] = 8'd6;
        rom[275][25] = 8'd24;
        rom[275][26] = -8'd21;
        rom[275][27] = -8'd43;
        rom[275][28] = 8'd23;
        rom[275][29] = -8'd11;
        rom[275][30] = -8'd27;
        rom[275][31] = 8'd9;
        rom[275][32] = -8'd28;
        rom[275][33] = -8'd21;
        rom[275][34] = 8'd14;
        rom[275][35] = 8'd4;
        rom[275][36] = 8'd4;
        rom[275][37] = 8'd7;
        rom[275][38] = -8'd24;
        rom[275][39] = -8'd31;
        rom[275][40] = -8'd16;
        rom[275][41] = -8'd10;
        rom[275][42] = -8'd13;
        rom[275][43] = -8'd71;
        rom[275][44] = 8'd16;
        rom[275][45] = -8'd4;
        rom[275][46] = 8'd3;
        rom[275][47] = 8'd29;
        rom[275][48] = -8'd11;
        rom[275][49] = 8'd2;
        rom[275][50] = -8'd5;
        rom[275][51] = 8'd21;
        rom[275][52] = -8'd1;
        rom[275][53] = 8'd6;
        rom[275][54] = -8'd34;
        rom[275][55] = -8'd37;
        rom[275][56] = -8'd31;
        rom[275][57] = 8'd7;
        rom[275][58] = 8'd22;
        rom[275][59] = 8'd2;
        rom[275][60] = -8'd2;
        rom[275][61] = -8'd5;
        rom[275][62] = 8'd3;
        rom[275][63] = -8'd26;
        rom[276][0] = -8'd4;
        rom[276][1] = 8'd5;
        rom[276][2] = -8'd24;
        rom[276][3] = 8'd13;
        rom[276][4] = -8'd22;
        rom[276][5] = -8'd5;
        rom[276][6] = -8'd18;
        rom[276][7] = -8'd35;
        rom[276][8] = 8'd3;
        rom[276][9] = 8'd10;
        rom[276][10] = -8'd4;
        rom[276][11] = -8'd10;
        rom[276][12] = -8'd6;
        rom[276][13] = -8'd17;
        rom[276][14] = -8'd35;
        rom[276][15] = -8'd25;
        rom[276][16] = -8'd18;
        rom[276][17] = 8'd10;
        rom[276][18] = -8'd45;
        rom[276][19] = 8'd9;
        rom[276][20] = -8'd2;
        rom[276][21] = -8'd2;
        rom[276][22] = -8'd27;
        rom[276][23] = -8'd24;
        rom[276][24] = 8'd7;
        rom[276][25] = -8'd57;
        rom[276][26] = 8'd0;
        rom[276][27] = 8'd5;
        rom[276][28] = -8'd17;
        rom[276][29] = 8'd22;
        rom[276][30] = -8'd51;
        rom[276][31] = -8'd19;
        rom[276][32] = -8'd50;
        rom[276][33] = 8'd3;
        rom[276][34] = -8'd28;
        rom[276][35] = -8'd71;
        rom[276][36] = -8'd60;
        rom[276][37] = 8'd9;
        rom[276][38] = -8'd9;
        rom[276][39] = -8'd9;
        rom[276][40] = -8'd9;
        rom[276][41] = 8'd12;
        rom[276][42] = 8'd14;
        rom[276][43] = -8'd7;
        rom[276][44] = -8'd1;
        rom[276][45] = -8'd9;
        rom[276][46] = 8'd1;
        rom[276][47] = -8'd3;
        rom[276][48] = -8'd40;
        rom[276][49] = 8'd8;
        rom[276][50] = -8'd9;
        rom[276][51] = 8'd10;
        rom[276][52] = -8'd41;
        rom[276][53] = -8'd24;
        rom[276][54] = -8'd3;
        rom[276][55] = 8'd12;
        rom[276][56] = -8'd16;
        rom[276][57] = 8'd5;
        rom[276][58] = -8'd11;
        rom[276][59] = 8'd7;
        rom[276][60] = -8'd26;
        rom[276][61] = -8'd24;
        rom[276][62] = 8'd9;
        rom[276][63] = -8'd48;
        rom[277][0] = 8'd9;
        rom[277][1] = -8'd7;
        rom[277][2] = -8'd3;
        rom[277][3] = -8'd5;
        rom[277][4] = -8'd5;
        rom[277][5] = -8'd9;
        rom[277][6] = 8'd2;
        rom[277][7] = -8'd9;
        rom[277][8] = -8'd7;
        rom[277][9] = 8'd3;
        rom[277][10] = -8'd2;
        rom[277][11] = -8'd5;
        rom[277][12] = -8'd8;
        rom[277][13] = 8'd3;
        rom[277][14] = 8'd2;
        rom[277][15] = -8'd1;
        rom[277][16] = -8'd2;
        rom[277][17] = 8'd6;
        rom[277][18] = 8'd5;
        rom[277][19] = -8'd7;
        rom[277][20] = 8'd2;
        rom[277][21] = -8'd5;
        rom[277][22] = -8'd3;
        rom[277][23] = 8'd4;
        rom[277][24] = 8'd6;
        rom[277][25] = 8'd7;
        rom[277][26] = -8'd9;
        rom[277][27] = 8'd0;
        rom[277][28] = -8'd8;
        rom[277][29] = -8'd3;
        rom[277][30] = -8'd1;
        rom[277][31] = 8'd1;
        rom[277][32] = 8'd3;
        rom[277][33] = -8'd9;
        rom[277][34] = 8'd1;
        rom[277][35] = 8'd10;
        rom[277][36] = 8'd4;
        rom[277][37] = 8'd8;
        rom[277][38] = 8'd5;
        rom[277][39] = 8'd9;
        rom[277][40] = 8'd4;
        rom[277][41] = 8'd5;
        rom[277][42] = -8'd2;
        rom[277][43] = 8'd4;
        rom[277][44] = -8'd3;
        rom[277][45] = 8'd8;
        rom[277][46] = -8'd1;
        rom[277][47] = -8'd1;
        rom[277][48] = 8'd1;
        rom[277][49] = 8'd5;
        rom[277][50] = 8'd10;
        rom[277][51] = -8'd2;
        rom[277][52] = -8'd3;
        rom[277][53] = 8'd2;
        rom[277][54] = 8'd9;
        rom[277][55] = 8'd5;
        rom[277][56] = -8'd3;
        rom[277][57] = -8'd11;
        rom[277][58] = 8'd1;
        rom[277][59] = -8'd8;
        rom[277][60] = 8'd6;
        rom[277][61] = -8'd9;
        rom[277][62] = -8'd6;
        rom[277][63] = 8'd12;
        rom[278][0] = -8'd39;
        rom[278][1] = 8'd17;
        rom[278][2] = 8'd0;
        rom[278][3] = -8'd31;
        rom[278][4] = -8'd48;
        rom[278][5] = -8'd36;
        rom[278][6] = -8'd19;
        rom[278][7] = 8'd26;
        rom[278][8] = 8'd8;
        rom[278][9] = -8'd18;
        rom[278][10] = 8'd13;
        rom[278][11] = 8'd8;
        rom[278][12] = -8'd24;
        rom[278][13] = 8'd13;
        rom[278][14] = 8'd8;
        rom[278][15] = -8'd29;
        rom[278][16] = 8'd36;
        rom[278][17] = 8'd15;
        rom[278][18] = -8'd46;
        rom[278][19] = 8'd8;
        rom[278][20] = -8'd3;
        rom[278][21] = -8'd7;
        rom[278][22] = 8'd33;
        rom[278][23] = -8'd43;
        rom[278][24] = -8'd3;
        rom[278][25] = 8'd21;
        rom[278][26] = -8'd9;
        rom[278][27] = 8'd14;
        rom[278][28] = -8'd5;
        rom[278][29] = -8'd22;
        rom[278][30] = -8'd15;
        rom[278][31] = -8'd23;
        rom[278][32] = -8'd11;
        rom[278][33] = 8'd37;
        rom[278][34] = 8'd13;
        rom[278][35] = -8'd18;
        rom[278][36] = 8'd11;
        rom[278][37] = 8'd30;
        rom[278][38] = 8'd33;
        rom[278][39] = -8'd9;
        rom[278][40] = -8'd6;
        rom[278][41] = -8'd15;
        rom[278][42] = 8'd17;
        rom[278][43] = -8'd15;
        rom[278][44] = -8'd49;
        rom[278][45] = 8'd7;
        rom[278][46] = 8'd19;
        rom[278][47] = -8'd111;
        rom[278][48] = -8'd35;
        rom[278][49] = -8'd40;
        rom[278][50] = -8'd36;
        rom[278][51] = 8'd18;
        rom[278][52] = 8'd10;
        rom[278][53] = -8'd38;
        rom[278][54] = -8'd23;
        rom[278][55] = -8'd17;
        rom[278][56] = -8'd34;
        rom[278][57] = 8'd14;
        rom[278][58] = -8'd21;
        rom[278][59] = 8'd19;
        rom[278][60] = -8'd31;
        rom[278][61] = -8'd5;
        rom[278][62] = -8'd31;
        rom[278][63] = -8'd12;
        rom[279][0] = -8'd4;
        rom[279][1] = 8'd4;
        rom[279][2] = -8'd19;
        rom[279][3] = -8'd15;
        rom[279][4] = 8'd25;
        rom[279][5] = 8'd12;
        rom[279][6] = 8'd8;
        rom[279][7] = -8'd12;
        rom[279][8] = 8'd5;
        rom[279][9] = -8'd1;
        rom[279][10] = -8'd14;
        rom[279][11] = 8'd2;
        rom[279][12] = 8'd40;
        rom[279][13] = 8'd38;
        rom[279][14] = -8'd29;
        rom[279][15] = -8'd36;
        rom[279][16] = -8'd8;
        rom[279][17] = -8'd18;
        rom[279][18] = -8'd15;
        rom[279][19] = 8'd11;
        rom[279][20] = -8'd3;
        rom[279][21] = 8'd11;
        rom[279][22] = 8'd11;
        rom[279][23] = -8'd9;
        rom[279][24] = -8'd4;
        rom[279][25] = -8'd40;
        rom[279][26] = -8'd19;
        rom[279][27] = 8'd8;
        rom[279][28] = 8'd36;
        rom[279][29] = 8'd25;
        rom[279][30] = -8'd12;
        rom[279][31] = 8'd10;
        rom[279][32] = -8'd7;
        rom[279][33] = 8'd1;
        rom[279][34] = -8'd14;
        rom[279][35] = -8'd27;
        rom[279][36] = -8'd4;
        rom[279][37] = -8'd14;
        rom[279][38] = 8'd30;
        rom[279][39] = -8'd6;
        rom[279][40] = -8'd3;
        rom[279][41] = 8'd13;
        rom[279][42] = -8'd7;
        rom[279][43] = -8'd11;
        rom[279][44] = -8'd27;
        rom[279][45] = -8'd14;
        rom[279][46] = -8'd2;
        rom[279][47] = 8'd42;
        rom[279][48] = -8'd62;
        rom[279][49] = -8'd12;
        rom[279][50] = -8'd23;
        rom[279][51] = -8'd16;
        rom[279][52] = -8'd7;
        rom[279][53] = 8'd1;
        rom[279][54] = 8'd24;
        rom[279][55] = -8'd2;
        rom[279][56] = 8'd27;
        rom[279][57] = -8'd11;
        rom[279][58] = 8'd17;
        rom[279][59] = -8'd11;
        rom[279][60] = -8'd22;
        rom[279][61] = 8'd0;
        rom[279][62] = -8'd47;
        rom[279][63] = 8'd17;
        rom[280][0] = 8'd19;
        rom[280][1] = 8'd12;
        rom[280][2] = -8'd6;
        rom[280][3] = 8'd26;
        rom[280][4] = -8'd22;
        rom[280][5] = 8'd2;
        rom[280][6] = 8'd3;
        rom[280][7] = 8'd26;
        rom[280][8] = -8'd12;
        rom[280][9] = -8'd6;
        rom[280][10] = -8'd19;
        rom[280][11] = 8'd1;
        rom[280][12] = 8'd31;
        rom[280][13] = 8'd27;
        rom[280][14] = -8'd27;
        rom[280][15] = 8'd17;
        rom[280][16] = -8'd3;
        rom[280][17] = 8'd3;
        rom[280][18] = -8'd5;
        rom[280][19] = 8'd33;
        rom[280][20] = -8'd4;
        rom[280][21] = 8'd6;
        rom[280][22] = -8'd33;
        rom[280][23] = 8'd47;
        rom[280][24] = -8'd31;
        rom[280][25] = -8'd10;
        rom[280][26] = 8'd12;
        rom[280][27] = 8'd23;
        rom[280][28] = 8'd18;
        rom[280][29] = 8'd2;
        rom[280][30] = 8'd8;
        rom[280][31] = -8'd4;
        rom[280][32] = 8'd3;
        rom[280][33] = 8'd25;
        rom[280][34] = -8'd9;
        rom[280][35] = -8'd5;
        rom[280][36] = -8'd7;
        rom[280][37] = 8'd38;
        rom[280][38] = -8'd14;
        rom[280][39] = -8'd3;
        rom[280][40] = 8'd7;
        rom[280][41] = 8'd5;
        rom[280][42] = 8'd3;
        rom[280][43] = 8'd15;
        rom[280][44] = -8'd20;
        rom[280][45] = 8'd8;
        rom[280][46] = 8'd15;
        rom[280][47] = -8'd18;
        rom[280][48] = -8'd1;
        rom[280][49] = 8'd7;
        rom[280][50] = -8'd6;
        rom[280][51] = -8'd7;
        rom[280][52] = 8'd3;
        rom[280][53] = -8'd4;
        rom[280][54] = -8'd1;
        rom[280][55] = 8'd12;
        rom[280][56] = 8'd13;
        rom[280][57] = -8'd15;
        rom[280][58] = -8'd30;
        rom[280][59] = -8'd2;
        rom[280][60] = -8'd20;
        rom[280][61] = 8'd2;
        rom[280][62] = -8'd17;
        rom[280][63] = 8'd2;
        rom[281][0] = 8'd24;
        rom[281][1] = 8'd4;
        rom[281][2] = -8'd48;
        rom[281][3] = 8'd0;
        rom[281][4] = -8'd86;
        rom[281][5] = -8'd3;
        rom[281][6] = 8'd22;
        rom[281][7] = -8'd7;
        rom[281][8] = -8'd3;
        rom[281][9] = -8'd3;
        rom[281][10] = -8'd33;
        rom[281][11] = 8'd14;
        rom[281][12] = 8'd29;
        rom[281][13] = -8'd33;
        rom[281][14] = -8'd11;
        rom[281][15] = 8'd20;
        rom[281][16] = 8'd13;
        rom[281][17] = 8'd23;
        rom[281][18] = 8'd16;
        rom[281][19] = -8'd15;
        rom[281][20] = 8'd0;
        rom[281][21] = -8'd40;
        rom[281][22] = 8'd13;
        rom[281][23] = 8'd19;
        rom[281][24] = -8'd14;
        rom[281][25] = 8'd44;
        rom[281][26] = 8'd47;
        rom[281][27] = -8'd29;
        rom[281][28] = 8'd8;
        rom[281][29] = 8'd19;
        rom[281][30] = -8'd3;
        rom[281][31] = 8'd34;
        rom[281][32] = 8'd24;
        rom[281][33] = 8'd2;
        rom[281][34] = -8'd47;
        rom[281][35] = -8'd16;
        rom[281][36] = 8'd46;
        rom[281][37] = 8'd22;
        rom[281][38] = 8'd18;
        rom[281][39] = -8'd10;
        rom[281][40] = -8'd46;
        rom[281][41] = -8'd10;
        rom[281][42] = 8'd0;
        rom[281][43] = -8'd20;
        rom[281][44] = 8'd3;
        rom[281][45] = 8'd11;
        rom[281][46] = 8'd22;
        rom[281][47] = -8'd48;
        rom[281][48] = 8'd1;
        rom[281][49] = -8'd2;
        rom[281][50] = -8'd52;
        rom[281][51] = -8'd10;
        rom[281][52] = -8'd36;
        rom[281][53] = -8'd36;
        rom[281][54] = -8'd11;
        rom[281][55] = -8'd12;
        rom[281][56] = -8'd5;
        rom[281][57] = -8'd40;
        rom[281][58] = 8'd32;
        rom[281][59] = 8'd26;
        rom[281][60] = 8'd26;
        rom[281][61] = -8'd13;
        rom[281][62] = 8'd0;
        rom[281][63] = 8'd12;
        rom[282][0] = -8'd6;
        rom[282][1] = -8'd7;
        rom[282][2] = 8'd23;
        rom[282][3] = -8'd51;
        rom[282][4] = 8'd9;
        rom[282][5] = 8'd26;
        rom[282][6] = 8'd35;
        rom[282][7] = -8'd39;
        rom[282][8] = 8'd16;
        rom[282][9] = 8'd8;
        rom[282][10] = 8'd27;
        rom[282][11] = -8'd47;
        rom[282][12] = -8'd52;
        rom[282][13] = 8'd5;
        rom[282][14] = 8'd23;
        rom[282][15] = -8'd66;
        rom[282][16] = 8'd3;
        rom[282][17] = 8'd15;
        rom[282][18] = 8'd2;
        rom[282][19] = 8'd5;
        rom[282][20] = -8'd12;
        rom[282][21] = 8'd6;
        rom[282][22] = 8'd10;
        rom[282][23] = -8'd26;
        rom[282][24] = -8'd16;
        rom[282][25] = 8'd15;
        rom[282][26] = 8'd19;
        rom[282][27] = -8'd42;
        rom[282][28] = -8'd4;
        rom[282][29] = -8'd4;
        rom[282][30] = -8'd13;
        rom[282][31] = -8'd20;
        rom[282][32] = 8'd6;
        rom[282][33] = 8'd22;
        rom[282][34] = 8'd4;
        rom[282][35] = 8'd19;
        rom[282][36] = 8'd6;
        rom[282][37] = 8'd4;
        rom[282][38] = 8'd13;
        rom[282][39] = 8'd0;
        rom[282][40] = 8'd27;
        rom[282][41] = 8'd16;
        rom[282][42] = 8'd3;
        rom[282][43] = -8'd7;
        rom[282][44] = 8'd13;
        rom[282][45] = -8'd46;
        rom[282][46] = 8'd3;
        rom[282][47] = 8'd0;
        rom[282][48] = -8'd6;
        rom[282][49] = -8'd13;
        rom[282][50] = -8'd6;
        rom[282][51] = -8'd20;
        rom[282][52] = -8'd32;
        rom[282][53] = -8'd14;
        rom[282][54] = -8'd52;
        rom[282][55] = -8'd29;
        rom[282][56] = -8'd1;
        rom[282][57] = -8'd23;
        rom[282][58] = -8'd27;
        rom[282][59] = 8'd2;
        rom[282][60] = 8'd23;
        rom[282][61] = 8'd0;
        rom[282][62] = -8'd8;
        rom[282][63] = -8'd20;
        rom[283][0] = -8'd5;
        rom[283][1] = -8'd21;
        rom[283][2] = 8'd20;
        rom[283][3] = -8'd16;
        rom[283][4] = 8'd11;
        rom[283][5] = 8'd52;
        rom[283][6] = -8'd16;
        rom[283][7] = 8'd3;
        rom[283][8] = 8'd33;
        rom[283][9] = 8'd22;
        rom[283][10] = -8'd50;
        rom[283][11] = -8'd21;
        rom[283][12] = -8'd65;
        rom[283][13] = 8'd3;
        rom[283][14] = 8'd0;
        rom[283][15] = 8'd8;
        rom[283][16] = -8'd7;
        rom[283][17] = 8'd8;
        rom[283][18] = 8'd28;
        rom[283][19] = -8'd18;
        rom[283][20] = -8'd10;
        rom[283][21] = -8'd32;
        rom[283][22] = 8'd14;
        rom[283][23] = 8'd6;
        rom[283][24] = 8'd6;
        rom[283][25] = 8'd36;
        rom[283][26] = 8'd16;
        rom[283][27] = 8'd0;
        rom[283][28] = 8'd4;
        rom[283][29] = 8'd10;
        rom[283][30] = 8'd6;
        rom[283][31] = -8'd25;
        rom[283][32] = 8'd24;
        rom[283][33] = 8'd19;
        rom[283][34] = -8'd63;
        rom[283][35] = 8'd25;
        rom[283][36] = -8'd2;
        rom[283][37] = 8'd22;
        rom[283][38] = 8'd10;
        rom[283][39] = -8'd20;
        rom[283][40] = 8'd5;
        rom[283][41] = -8'd23;
        rom[283][42] = 8'd3;
        rom[283][43] = -8'd44;
        rom[283][44] = -8'd45;
        rom[283][45] = 8'd41;
        rom[283][46] = 8'd53;
        rom[283][47] = -8'd38;
        rom[283][48] = -8'd45;
        rom[283][49] = -8'd18;
        rom[283][50] = 8'd4;
        rom[283][51] = 8'd31;
        rom[283][52] = 8'd7;
        rom[283][53] = 8'd5;
        rom[283][54] = -8'd4;
        rom[283][55] = 8'd23;
        rom[283][56] = -8'd6;
        rom[283][57] = -8'd39;
        rom[283][58] = 8'd12;
        rom[283][59] = 8'd38;
        rom[283][60] = 8'd10;
        rom[283][61] = -8'd26;
        rom[283][62] = 8'd12;
        rom[283][63] = -8'd34;
        rom[284][0] = -8'd78;
        rom[284][1] = -8'd17;
        rom[284][2] = -8'd36;
        rom[284][3] = -8'd36;
        rom[284][4] = -8'd5;
        rom[284][5] = -8'd37;
        rom[284][6] = -8'd4;
        rom[284][7] = 8'd32;
        rom[284][8] = -8'd7;
        rom[284][9] = 8'd16;
        rom[284][10] = 8'd23;
        rom[284][11] = -8'd14;
        rom[284][12] = -8'd55;
        rom[284][13] = -8'd33;
        rom[284][14] = -8'd22;
        rom[284][15] = 8'd18;
        rom[284][16] = -8'd11;
        rom[284][17] = -8'd5;
        rom[284][18] = -8'd21;
        rom[284][19] = -8'd70;
        rom[284][20] = -8'd9;
        rom[284][21] = -8'd42;
        rom[284][22] = -8'd31;
        rom[284][23] = -8'd12;
        rom[284][24] = -8'd25;
        rom[284][25] = 8'd20;
        rom[284][26] = -8'd52;
        rom[284][27] = -8'd31;
        rom[284][28] = -8'd14;
        rom[284][29] = 8'd15;
        rom[284][30] = 8'd15;
        rom[284][31] = 8'd1;
        rom[284][32] = -8'd37;
        rom[284][33] = -8'd54;
        rom[284][34] = 8'd17;
        rom[284][35] = 8'd8;
        rom[284][36] = 8'd11;
        rom[284][37] = 8'd2;
        rom[284][38] = -8'd2;
        rom[284][39] = -8'd11;
        rom[284][40] = -8'd40;
        rom[284][41] = -8'd4;
        rom[284][42] = -8'd24;
        rom[284][43] = -8'd27;
        rom[284][44] = 8'd26;
        rom[284][45] = 8'd13;
        rom[284][46] = -8'd8;
        rom[284][47] = -8'd1;
        rom[284][48] = -8'd22;
        rom[284][49] = 8'd1;
        rom[284][50] = -8'd7;
        rom[284][51] = 8'd14;
        rom[284][52] = -8'd5;
        rom[284][53] = -8'd8;
        rom[284][54] = -8'd42;
        rom[284][55] = -8'd24;
        rom[284][56] = 8'd7;
        rom[284][57] = 8'd1;
        rom[284][58] = 8'd6;
        rom[284][59] = -8'd5;
        rom[284][60] = 8'd22;
        rom[284][61] = 8'd24;
        rom[284][62] = 8'd10;
        rom[284][63] = -8'd13;
        rom[285][0] = 8'd13;
        rom[285][1] = -8'd67;
        rom[285][2] = -8'd15;
        rom[285][3] = -8'd20;
        rom[285][4] = 8'd28;
        rom[285][5] = -8'd5;
        rom[285][6] = -8'd5;
        rom[285][7] = -8'd1;
        rom[285][8] = 8'd20;
        rom[285][9] = -8'd3;
        rom[285][10] = 8'd42;
        rom[285][11] = 8'd5;
        rom[285][12] = -8'd22;
        rom[285][13] = 8'd45;
        rom[285][14] = 8'd14;
        rom[285][15] = -8'd28;
        rom[285][16] = 8'd30;
        rom[285][17] = 8'd2;
        rom[285][18] = -8'd5;
        rom[285][19] = -8'd49;
        rom[285][20] = -8'd12;
        rom[285][21] = 8'd6;
        rom[285][22] = -8'd17;
        rom[285][23] = 8'd1;
        rom[285][24] = -8'd49;
        rom[285][25] = 8'd10;
        rom[285][26] = 8'd5;
        rom[285][27] = -8'd81;
        rom[285][28] = -8'd5;
        rom[285][29] = -8'd16;
        rom[285][30] = -8'd25;
        rom[285][31] = -8'd17;
        rom[285][32] = -8'd15;
        rom[285][33] = 8'd18;
        rom[285][34] = -8'd8;
        rom[285][35] = -8'd9;
        rom[285][36] = -8'd4;
        rom[285][37] = -8'd2;
        rom[285][38] = -8'd89;
        rom[285][39] = -8'd14;
        rom[285][40] = -8'd20;
        rom[285][41] = -8'd26;
        rom[285][42] = -8'd19;
        rom[285][43] = -8'd15;
        rom[285][44] = -8'd2;
        rom[285][45] = 8'd23;
        rom[285][46] = 8'd10;
        rom[285][47] = 8'd36;
        rom[285][48] = -8'd27;
        rom[285][49] = -8'd20;
        rom[285][50] = 8'd0;
        rom[285][51] = 8'd24;
        rom[285][52] = 8'd6;
        rom[285][53] = -8'd22;
        rom[285][54] = -8'd50;
        rom[285][55] = 8'd4;
        rom[285][56] = -8'd46;
        rom[285][57] = -8'd3;
        rom[285][58] = 8'd0;
        rom[285][59] = -8'd30;
        rom[285][60] = -8'd68;
        rom[285][61] = 8'd10;
        rom[285][62] = -8'd20;
        rom[285][63] = -8'd13;
        rom[286][0] = 8'd6;
        rom[286][1] = -8'd31;
        rom[286][2] = -8'd5;
        rom[286][3] = 8'd15;
        rom[286][4] = 8'd13;
        rom[286][5] = 8'd24;
        rom[286][6] = 8'd16;
        rom[286][7] = -8'd11;
        rom[286][8] = -8'd2;
        rom[286][9] = 8'd2;
        rom[286][10] = 8'd19;
        rom[286][11] = 8'd29;
        rom[286][12] = 8'd5;
        rom[286][13] = 8'd5;
        rom[286][14] = -8'd19;
        rom[286][15] = -8'd11;
        rom[286][16] = -8'd4;
        rom[286][17] = 8'd42;
        rom[286][18] = 8'd10;
        rom[286][19] = -8'd3;
        rom[286][20] = -8'd6;
        rom[286][21] = 8'd0;
        rom[286][22] = 8'd5;
        rom[286][23] = 8'd7;
        rom[286][24] = -8'd21;
        rom[286][25] = -8'd53;
        rom[286][26] = 8'd10;
        rom[286][27] = -8'd48;
        rom[286][28] = 8'd7;
        rom[286][29] = 8'd14;
        rom[286][30] = 8'd23;
        rom[286][31] = -8'd25;
        rom[286][32] = 8'd4;
        rom[286][33] = -8'd31;
        rom[286][34] = -8'd35;
        rom[286][35] = -8'd18;
        rom[286][36] = 8'd5;
        rom[286][37] = -8'd1;
        rom[286][38] = 8'd21;
        rom[286][39] = 8'd2;
        rom[286][40] = -8'd37;
        rom[286][41] = -8'd3;
        rom[286][42] = 8'd8;
        rom[286][43] = -8'd65;
        rom[286][44] = 8'd13;
        rom[286][45] = 8'd7;
        rom[286][46] = 8'd1;
        rom[286][47] = 8'd12;
        rom[286][48] = -8'd27;
        rom[286][49] = -8'd20;
        rom[286][50] = -8'd15;
        rom[286][51] = -8'd44;
        rom[286][52] = -8'd1;
        rom[286][53] = -8'd25;
        rom[286][54] = -8'd59;
        rom[286][55] = -8'd19;
        rom[286][56] = -8'd31;
        rom[286][57] = 8'd1;
        rom[286][58] = 8'd21;
        rom[286][59] = 8'd7;
        rom[286][60] = 8'd23;
        rom[286][61] = 8'd10;
        rom[286][62] = 8'd20;
        rom[286][63] = 8'd7;
        rom[287][0] = 8'd9;
        rom[287][1] = -8'd22;
        rom[287][2] = -8'd22;
        rom[287][3] = -8'd28;
        rom[287][4] = -8'd11;
        rom[287][5] = -8'd22;
        rom[287][6] = -8'd32;
        rom[287][7] = 8'd4;
        rom[287][8] = -8'd34;
        rom[287][9] = -8'd9;
        rom[287][10] = -8'd5;
        rom[287][11] = -8'd49;
        rom[287][12] = 8'd10;
        rom[287][13] = -8'd31;
        rom[287][14] = 8'd30;
        rom[287][15] = 8'd25;
        rom[287][16] = 8'd30;
        rom[287][17] = 8'd25;
        rom[287][18] = -8'd42;
        rom[287][19] = 8'd3;
        rom[287][20] = -8'd7;
        rom[287][21] = -8'd36;
        rom[287][22] = -8'd13;
        rom[287][23] = -8'd22;
        rom[287][24] = -8'd14;
        rom[287][25] = 8'd25;
        rom[287][26] = 8'd5;
        rom[287][27] = -8'd39;
        rom[287][28] = 8'd19;
        rom[287][29] = -8'd32;
        rom[287][30] = 8'd23;
        rom[287][31] = 8'd2;
        rom[287][32] = -8'd21;
        rom[287][33] = 8'd12;
        rom[287][34] = 8'd3;
        rom[287][35] = -8'd25;
        rom[287][36] = 8'd1;
        rom[287][37] = 8'd34;
        rom[287][38] = -8'd4;
        rom[287][39] = 8'd14;
        rom[287][40] = 8'd0;
        rom[287][41] = 8'd1;
        rom[287][42] = 8'd11;
        rom[287][43] = -8'd9;
        rom[287][44] = -8'd28;
        rom[287][45] = -8'd50;
        rom[287][46] = -8'd8;
        rom[287][47] = -8'd33;
        rom[287][48] = 8'd32;
        rom[287][49] = 8'd13;
        rom[287][50] = 8'd7;
        rom[287][51] = -8'd31;
        rom[287][52] = -8'd12;
        rom[287][53] = 8'd3;
        rom[287][54] = -8'd60;
        rom[287][55] = -8'd39;
        rom[287][56] = -8'd26;
        rom[287][57] = 8'd17;
        rom[287][58] = -8'd16;
        rom[287][59] = -8'd17;
        rom[287][60] = -8'd24;
        rom[287][61] = -8'd4;
        rom[287][62] = -8'd11;
        rom[287][63] = 8'd40;
        rom[288][0] = 8'd32;
        rom[288][1] = -8'd4;
        rom[288][2] = 8'd21;
        rom[288][3] = 8'd17;
        rom[288][4] = -8'd16;
        rom[288][5] = 8'd23;
        rom[288][6] = 8'd23;
        rom[288][7] = 8'd29;
        rom[288][8] = 8'd11;
        rom[288][9] = 8'd25;
        rom[288][10] = -8'd35;
        rom[288][11] = -8'd5;
        rom[288][12] = -8'd15;
        rom[288][13] = -8'd43;
        rom[288][14] = 8'd10;
        rom[288][15] = -8'd31;
        rom[288][16] = -8'd27;
        rom[288][17] = 8'd7;
        rom[288][18] = 8'd7;
        rom[288][19] = 8'd13;
        rom[288][20] = -8'd11;
        rom[288][21] = -8'd7;
        rom[288][22] = -8'd20;
        rom[288][23] = -8'd4;
        rom[288][24] = 8'd22;
        rom[288][25] = -8'd27;
        rom[288][26] = 8'd3;
        rom[288][27] = -8'd31;
        rom[288][28] = -8'd10;
        rom[288][29] = 8'd2;
        rom[288][30] = -8'd20;
        rom[288][31] = -8'd22;
        rom[288][32] = 8'd16;
        rom[288][33] = -8'd35;
        rom[288][34] = -8'd59;
        rom[288][35] = 8'd3;
        rom[288][36] = -8'd16;
        rom[288][37] = -8'd43;
        rom[288][38] = -8'd10;
        rom[288][39] = -8'd30;
        rom[288][40] = 8'd23;
        rom[288][41] = -8'd22;
        rom[288][42] = -8'd17;
        rom[288][43] = -8'd8;
        rom[288][44] = -8'd12;
        rom[288][45] = 8'd20;
        rom[288][46] = -8'd18;
        rom[288][47] = -8'd50;
        rom[288][48] = -8'd23;
        rom[288][49] = 8'd23;
        rom[288][50] = 8'd28;
        rom[288][51] = 8'd28;
        rom[288][52] = 8'd2;
        rom[288][53] = -8'd1;
        rom[288][54] = 8'd4;
        rom[288][55] = 8'd11;
        rom[288][56] = 8'd7;
        rom[288][57] = 8'd7;
        rom[288][58] = -8'd12;
        rom[288][59] = 8'd20;
        rom[288][60] = 8'd35;
        rom[288][61] = -8'd10;
        rom[288][62] = 8'd10;
        rom[288][63] = 8'd29;
        rom[289][0] = 8'd3;
        rom[289][1] = -8'd31;
        rom[289][2] = 8'd4;
        rom[289][3] = -8'd10;
        rom[289][4] = -8'd14;
        rom[289][5] = -8'd7;
        rom[289][6] = -8'd30;
        rom[289][7] = 8'd6;
        rom[289][8] = 8'd3;
        rom[289][9] = -8'd15;
        rom[289][10] = 8'd27;
        rom[289][11] = 8'd4;
        rom[289][12] = 8'd7;
        rom[289][13] = -8'd18;
        rom[289][14] = -8'd9;
        rom[289][15] = 8'd29;
        rom[289][16] = 8'd29;
        rom[289][17] = 8'd28;
        rom[289][18] = 8'd3;
        rom[289][19] = -8'd19;
        rom[289][20] = -8'd8;
        rom[289][21] = 8'd6;
        rom[289][22] = -8'd10;
        rom[289][23] = -8'd17;
        rom[289][24] = -8'd34;
        rom[289][25] = 8'd31;
        rom[289][26] = -8'd19;
        rom[289][27] = 8'd10;
        rom[289][28] = 8'd14;
        rom[289][29] = 8'd44;
        rom[289][30] = 8'd16;
        rom[289][31] = -8'd22;
        rom[289][32] = 8'd50;
        rom[289][33] = 8'd40;
        rom[289][34] = -8'd11;
        rom[289][35] = 8'd41;
        rom[289][36] = -8'd10;
        rom[289][37] = 8'd34;
        rom[289][38] = 8'd1;
        rom[289][39] = -8'd13;
        rom[289][40] = -8'd21;
        rom[289][41] = -8'd17;
        rom[289][42] = 8'd8;
        rom[289][43] = -8'd3;
        rom[289][44] = 8'd12;
        rom[289][45] = 8'd7;
        rom[289][46] = 8'd23;
        rom[289][47] = 8'd4;
        rom[289][48] = -8'd63;
        rom[289][49] = 8'd11;
        rom[289][50] = 8'd26;
        rom[289][51] = 8'd16;
        rom[289][52] = -8'd73;
        rom[289][53] = -8'd5;
        rom[289][54] = -8'd17;
        rom[289][55] = 8'd43;
        rom[289][56] = 8'd1;
        rom[289][57] = -8'd19;
        rom[289][58] = 8'd5;
        rom[289][59] = 8'd28;
        rom[289][60] = -8'd65;
        rom[289][61] = -8'd1;
        rom[289][62] = 8'd36;
        rom[289][63] = -8'd6;
        rom[290][0] = -8'd13;
        rom[290][1] = 8'd0;
        rom[290][2] = -8'd25;
        rom[290][3] = -8'd19;
        rom[290][4] = 8'd8;
        rom[290][5] = 8'd5;
        rom[290][6] = -8'd3;
        rom[290][7] = 8'd3;
        rom[290][8] = -8'd52;
        rom[290][9] = -8'd13;
        rom[290][10] = -8'd22;
        rom[290][11] = 8'd15;
        rom[290][12] = 8'd21;
        rom[290][13] = -8'd2;
        rom[290][14] = 8'd8;
        rom[290][15] = 8'd12;
        rom[290][16] = -8'd8;
        rom[290][17] = 8'd16;
        rom[290][18] = -8'd17;
        rom[290][19] = -8'd6;
        rom[290][20] = -8'd20;
        rom[290][21] = 8'd3;
        rom[290][22] = 8'd30;
        rom[290][23] = 8'd0;
        rom[290][24] = 8'd26;
        rom[290][25] = 8'd6;
        rom[290][26] = 8'd11;
        rom[290][27] = -8'd22;
        rom[290][28] = -8'd42;
        rom[290][29] = -8'd10;
        rom[290][30] = -8'd2;
        rom[290][31] = -8'd40;
        rom[290][32] = -8'd9;
        rom[290][33] = -8'd20;
        rom[290][34] = 8'd20;
        rom[290][35] = -8'd26;
        rom[290][36] = -8'd8;
        rom[290][37] = -8'd4;
        rom[290][38] = -8'd8;
        rom[290][39] = 8'd17;
        rom[290][40] = -8'd22;
        rom[290][41] = -8'd31;
        rom[290][42] = -8'd25;
        rom[290][43] = 8'd10;
        rom[290][44] = -8'd37;
        rom[290][45] = -8'd20;
        rom[290][46] = -8'd24;
        rom[290][47] = -8'd7;
        rom[290][48] = -8'd15;
        rom[290][49] = 8'd26;
        rom[290][50] = -8'd21;
        rom[290][51] = -8'd4;
        rom[290][52] = -8'd5;
        rom[290][53] = 8'd4;
        rom[290][54] = 8'd8;
        rom[290][55] = -8'd21;
        rom[290][56] = -8'd16;
        rom[290][57] = 8'd0;
        rom[290][58] = -8'd11;
        rom[290][59] = 8'd23;
        rom[290][60] = -8'd2;
        rom[290][61] = 8'd4;
        rom[290][62] = -8'd1;
        rom[290][63] = 8'd13;
        rom[291][0] = -8'd54;
        rom[291][1] = 8'd6;
        rom[291][2] = 8'd29;
        rom[291][3] = -8'd10;
        rom[291][4] = 8'd22;
        rom[291][5] = -8'd17;
        rom[291][6] = -8'd32;
        rom[291][7] = 8'd5;
        rom[291][8] = 8'd10;
        rom[291][9] = -8'd12;
        rom[291][10] = -8'd54;
        rom[291][11] = 8'd6;
        rom[291][12] = 8'd24;
        rom[291][13] = -8'd16;
        rom[291][14] = 8'd40;
        rom[291][15] = -8'd24;
        rom[291][16] = 8'd35;
        rom[291][17] = 8'd17;
        rom[291][18] = -8'd42;
        rom[291][19] = -8'd56;
        rom[291][20] = -8'd16;
        rom[291][21] = -8'd15;
        rom[291][22] = -8'd15;
        rom[291][23] = 8'd4;
        rom[291][24] = -8'd21;
        rom[291][25] = -8'd29;
        rom[291][26] = -8'd44;
        rom[291][27] = 8'd54;
        rom[291][28] = -8'd1;
        rom[291][29] = -8'd27;
        rom[291][30] = 8'd7;
        rom[291][31] = -8'd4;
        rom[291][32] = -8'd36;
        rom[291][33] = 8'd1;
        rom[291][34] = 8'd17;
        rom[291][35] = 8'd1;
        rom[291][36] = -8'd24;
        rom[291][37] = 8'd6;
        rom[291][38] = -8'd44;
        rom[291][39] = -8'd24;
        rom[291][40] = -8'd54;
        rom[291][41] = 8'd1;
        rom[291][42] = -8'd38;
        rom[291][43] = 8'd10;
        rom[291][44] = -8'd28;
        rom[291][45] = -8'd14;
        rom[291][46] = 8'd4;
        rom[291][47] = 8'd7;
        rom[291][48] = -8'd18;
        rom[291][49] = 8'd18;
        rom[291][50] = -8'd7;
        rom[291][51] = -8'd4;
        rom[291][52] = -8'd33;
        rom[291][53] = -8'd47;
        rom[291][54] = -8'd7;
        rom[291][55] = -8'd37;
        rom[291][56] = 8'd7;
        rom[291][57] = 8'd5;
        rom[291][58] = 8'd9;
        rom[291][59] = 8'd12;
        rom[291][60] = -8'd82;
        rom[291][61] = -8'd22;
        rom[291][62] = -8'd6;
        rom[291][63] = -8'd3;
        rom[292][0] = -8'd31;
        rom[292][1] = -8'd37;
        rom[292][2] = 8'd7;
        rom[292][3] = -8'd10;
        rom[292][4] = 8'd10;
        rom[292][5] = -8'd25;
        rom[292][6] = -8'd12;
        rom[292][7] = -8'd40;
        rom[292][8] = -8'd50;
        rom[292][9] = -8'd17;
        rom[292][10] = -8'd7;
        rom[292][11] = -8'd31;
        rom[292][12] = -8'd28;
        rom[292][13] = -8'd37;
        rom[292][14] = -8'd40;
        rom[292][15] = 8'd6;
        rom[292][16] = 8'd4;
        rom[292][17] = 8'd16;
        rom[292][18] = -8'd19;
        rom[292][19] = -8'd19;
        rom[292][20] = -8'd15;
        rom[292][21] = 8'd10;
        rom[292][22] = -8'd16;
        rom[292][23] = -8'd31;
        rom[292][24] = 8'd15;
        rom[292][25] = -8'd8;
        rom[292][26] = 8'd21;
        rom[292][27] = 8'd7;
        rom[292][28] = -8'd17;
        rom[292][29] = -8'd3;
        rom[292][30] = -8'd10;
        rom[292][31] = -8'd13;
        rom[292][32] = -8'd35;
        rom[292][33] = -8'd2;
        rom[292][34] = -8'd10;
        rom[292][35] = -8'd43;
        rom[292][36] = 8'd19;
        rom[292][37] = 8'd21;
        rom[292][38] = -8'd30;
        rom[292][39] = -8'd13;
        rom[292][40] = 8'd12;
        rom[292][41] = -8'd59;
        rom[292][42] = -8'd39;
        rom[292][43] = 8'd21;
        rom[292][44] = -8'd6;
        rom[292][45] = -8'd23;
        rom[292][46] = -8'd82;
        rom[292][47] = -8'd10;
        rom[292][48] = 8'd20;
        rom[292][49] = -8'd21;
        rom[292][50] = -8'd35;
        rom[292][51] = -8'd15;
        rom[292][52] = -8'd60;
        rom[292][53] = -8'd26;
        rom[292][54] = -8'd26;
        rom[292][55] = 8'd12;
        rom[292][56] = -8'd8;
        rom[292][57] = 8'd2;
        rom[292][58] = -8'd14;
        rom[292][59] = -8'd22;
        rom[292][60] = -8'd24;
        rom[292][61] = -8'd23;
        rom[292][62] = -8'd9;
        rom[292][63] = -8'd10;
        rom[293][0] = -8'd59;
        rom[293][1] = -8'd113;
        rom[293][2] = -8'd20;
        rom[293][3] = -8'd6;
        rom[293][4] = -8'd57;
        rom[293][5] = 8'd24;
        rom[293][6] = 8'd0;
        rom[293][7] = 8'd22;
        rom[293][8] = 8'd9;
        rom[293][9] = 8'd9;
        rom[293][10] = 8'd16;
        rom[293][11] = -8'd25;
        rom[293][12] = -8'd25;
        rom[293][13] = 8'd15;
        rom[293][14] = -8'd37;
        rom[293][15] = -8'd25;
        rom[293][16] = -8'd51;
        rom[293][17] = 8'd18;
        rom[293][18] = 8'd11;
        rom[293][19] = -8'd56;
        rom[293][20] = -8'd5;
        rom[293][21] = -8'd17;
        rom[293][22] = -8'd23;
        rom[293][23] = 8'd10;
        rom[293][24] = -8'd27;
        rom[293][25] = 8'd39;
        rom[293][26] = 8'd4;
        rom[293][27] = -8'd17;
        rom[293][28] = -8'd19;
        rom[293][29] = 8'd18;
        rom[293][30] = -8'd2;
        rom[293][31] = 8'd30;
        rom[293][32] = -8'd62;
        rom[293][33] = 8'd1;
        rom[293][34] = -8'd29;
        rom[293][35] = 8'd31;
        rom[293][36] = 8'd0;
        rom[293][37] = -8'd15;
        rom[293][38] = 8'd20;
        rom[293][39] = 8'd0;
        rom[293][40] = -8'd13;
        rom[293][41] = -8'd19;
        rom[293][42] = 8'd1;
        rom[293][43] = -8'd33;
        rom[293][44] = 8'd5;
        rom[293][45] = -8'd41;
        rom[293][46] = -8'd11;
        rom[293][47] = -8'd2;
        rom[293][48] = -8'd12;
        rom[293][49] = -8'd31;
        rom[293][50] = 8'd3;
        rom[293][51] = 8'd2;
        rom[293][52] = 8'd21;
        rom[293][53] = 8'd36;
        rom[293][54] = 8'd2;
        rom[293][55] = 8'd12;
        rom[293][56] = -8'd105;
        rom[293][57] = 8'd3;
        rom[293][58] = -8'd8;
        rom[293][59] = 8'd33;
        rom[293][60] = -8'd12;
        rom[293][61] = 8'd12;
        rom[293][62] = 8'd15;
        rom[293][63] = -8'd54;
        rom[294][0] = 8'd4;
        rom[294][1] = -8'd41;
        rom[294][2] = -8'd20;
        rom[294][3] = -8'd56;
        rom[294][4] = -8'd19;
        rom[294][5] = -8'd33;
        rom[294][6] = -8'd10;
        rom[294][7] = 8'd29;
        rom[294][8] = 8'd3;
        rom[294][9] = -8'd1;
        rom[294][10] = -8'd4;
        rom[294][11] = 8'd0;
        rom[294][12] = -8'd24;
        rom[294][13] = 8'd24;
        rom[294][14] = -8'd15;
        rom[294][15] = -8'd1;
        rom[294][16] = 8'd1;
        rom[294][17] = -8'd26;
        rom[294][18] = -8'd14;
        rom[294][19] = -8'd39;
        rom[294][20] = -8'd14;
        rom[294][21] = -8'd6;
        rom[294][22] = -8'd20;
        rom[294][23] = 8'd20;
        rom[294][24] = -8'd2;
        rom[294][25] = 8'd12;
        rom[294][26] = 8'd40;
        rom[294][27] = -8'd60;
        rom[294][28] = 8'd33;
        rom[294][29] = -8'd30;
        rom[294][30] = 8'd33;
        rom[294][31] = -8'd35;
        rom[294][32] = -8'd35;
        rom[294][33] = 8'd11;
        rom[294][34] = -8'd36;
        rom[294][35] = 8'd29;
        rom[294][36] = 8'd17;
        rom[294][37] = 8'd7;
        rom[294][38] = -8'd22;
        rom[294][39] = -8'd66;
        rom[294][40] = 8'd16;
        rom[294][41] = -8'd12;
        rom[294][42] = -8'd44;
        rom[294][43] = -8'd8;
        rom[294][44] = -8'd10;
        rom[294][45] = -8'd12;
        rom[294][46] = -8'd32;
        rom[294][47] = 8'd31;
        rom[294][48] = 8'd11;
        rom[294][49] = -8'd20;
        rom[294][50] = 8'd8;
        rom[294][51] = -8'd26;
        rom[294][52] = 8'd31;
        rom[294][53] = -8'd39;
        rom[294][54] = 8'd2;
        rom[294][55] = -8'd78;
        rom[294][56] = -8'd36;
        rom[294][57] = 8'd14;
        rom[294][58] = 8'd13;
        rom[294][59] = 8'd23;
        rom[294][60] = 8'd41;
        rom[294][61] = 8'd15;
        rom[294][62] = -8'd5;
        rom[294][63] = -8'd15;
        rom[295][0] = -8'd26;
        rom[295][1] = -8'd7;
        rom[295][2] = 8'd5;
        rom[295][3] = -8'd41;
        rom[295][4] = -8'd1;
        rom[295][5] = -8'd7;
        rom[295][6] = 8'd17;
        rom[295][7] = -8'd20;
        rom[295][8] = -8'd4;
        rom[295][9] = -8'd13;
        rom[295][10] = -8'd38;
        rom[295][11] = 8'd8;
        rom[295][12] = -8'd8;
        rom[295][13] = 8'd17;
        rom[295][14] = -8'd14;
        rom[295][15] = 8'd1;
        rom[295][16] = -8'd4;
        rom[295][17] = -8'd70;
        rom[295][18] = -8'd26;
        rom[295][19] = -8'd1;
        rom[295][20] = -8'd13;
        rom[295][21] = -8'd22;
        rom[295][22] = -8'd22;
        rom[295][23] = 8'd38;
        rom[295][24] = -8'd5;
        rom[295][25] = -8'd63;
        rom[295][26] = 8'd30;
        rom[295][27] = 8'd32;
        rom[295][28] = -8'd31;
        rom[295][29] = -8'd61;
        rom[295][30] = -8'd17;
        rom[295][31] = 8'd1;
        rom[295][32] = -8'd40;
        rom[295][33] = 8'd24;
        rom[295][34] = -8'd12;
        rom[295][35] = -8'd14;
        rom[295][36] = -8'd30;
        rom[295][37] = 8'd19;
        rom[295][38] = -8'd13;
        rom[295][39] = -8'd14;
        rom[295][40] = 8'd14;
        rom[295][41] = -8'd2;
        rom[295][42] = 8'd27;
        rom[295][43] = -8'd43;
        rom[295][44] = -8'd34;
        rom[295][45] = -8'd13;
        rom[295][46] = 8'd0;
        rom[295][47] = -8'd57;
        rom[295][48] = -8'd33;
        rom[295][49] = 8'd6;
        rom[295][50] = 8'd15;
        rom[295][51] = -8'd21;
        rom[295][52] = -8'd27;
        rom[295][53] = -8'd47;
        rom[295][54] = 8'd17;
        rom[295][55] = -8'd18;
        rom[295][56] = 8'd1;
        rom[295][57] = 8'd15;
        rom[295][58] = -8'd18;
        rom[295][59] = -8'd10;
        rom[295][60] = 8'd4;
        rom[295][61] = -8'd24;
        rom[295][62] = 8'd8;
        rom[295][63] = 8'd12;
        rom[296][0] = -8'd20;
        rom[296][1] = 8'd19;
        rom[296][2] = -8'd2;
        rom[296][3] = 8'd33;
        rom[296][4] = 8'd23;
        rom[296][5] = -8'd10;
        rom[296][6] = 8'd17;
        rom[296][7] = -8'd14;
        rom[296][8] = -8'd31;
        rom[296][9] = -8'd61;
        rom[296][10] = -8'd35;
        rom[296][11] = 8'd15;
        rom[296][12] = -8'd25;
        rom[296][13] = 8'd13;
        rom[296][14] = 8'd13;
        rom[296][15] = -8'd46;
        rom[296][16] = -8'd2;
        rom[296][17] = -8'd5;
        rom[296][18] = 8'd23;
        rom[296][19] = -8'd41;
        rom[296][20] = -8'd7;
        rom[296][21] = -8'd10;
        rom[296][22] = 8'd27;
        rom[296][23] = 8'd36;
        rom[296][24] = -8'd7;
        rom[296][25] = -8'd23;
        rom[296][26] = -8'd3;
        rom[296][27] = -8'd70;
        rom[296][28] = -8'd44;
        rom[296][29] = -8'd20;
        rom[296][30] = -8'd16;
        rom[296][31] = 8'd10;
        rom[296][32] = 8'd1;
        rom[296][33] = -8'd18;
        rom[296][34] = -8'd13;
        rom[296][35] = -8'd13;
        rom[296][36] = 8'd6;
        rom[296][37] = 8'd5;
        rom[296][38] = 8'd20;
        rom[296][39] = -8'd4;
        rom[296][40] = 8'd8;
        rom[296][41] = -8'd20;
        rom[296][42] = 8'd2;
        rom[296][43] = -8'd40;
        rom[296][44] = 8'd23;
        rom[296][45] = -8'd3;
        rom[296][46] = -8'd27;
        rom[296][47] = 8'd20;
        rom[296][48] = 8'd17;
        rom[296][49] = -8'd4;
        rom[296][50] = 8'd7;
        rom[296][51] = -8'd9;
        rom[296][52] = -8'd23;
        rom[296][53] = -8'd7;
        rom[296][54] = 8'd15;
        rom[296][55] = -8'd5;
        rom[296][56] = 8'd48;
        rom[296][57] = 8'd10;
        rom[296][58] = 8'd26;
        rom[296][59] = -8'd61;
        rom[296][60] = 8'd9;
        rom[296][61] = 8'd9;
        rom[296][62] = -8'd65;
        rom[296][63] = -8'd8;
        rom[297][0] = 8'd4;
        rom[297][1] = -8'd3;
        rom[297][2] = 8'd5;
        rom[297][3] = 8'd4;
        rom[297][4] = -8'd36;
        rom[297][5] = -8'd28;
        rom[297][6] = 8'd31;
        rom[297][7] = -8'd60;
        rom[297][8] = -8'd12;
        rom[297][9] = 8'd8;
        rom[297][10] = -8'd23;
        rom[297][11] = -8'd93;
        rom[297][12] = -8'd25;
        rom[297][13] = -8'd2;
        rom[297][14] = -8'd27;
        rom[297][15] = -8'd59;
        rom[297][16] = -8'd26;
        rom[297][17] = 8'd4;
        rom[297][18] = 8'd28;
        rom[297][19] = -8'd32;
        rom[297][20] = -8'd3;
        rom[297][21] = -8'd14;
        rom[297][22] = 8'd14;
        rom[297][23] = -8'd19;
        rom[297][24] = -8'd24;
        rom[297][25] = 8'd32;
        rom[297][26] = -8'd4;
        rom[297][27] = 8'd40;
        rom[297][28] = 8'd22;
        rom[297][29] = 8'd21;
        rom[297][30] = -8'd10;
        rom[297][31] = 8'd10;
        rom[297][32] = -8'd21;
        rom[297][33] = 8'd24;
        rom[297][34] = -8'd13;
        rom[297][35] = -8'd36;
        rom[297][36] = 8'd22;
        rom[297][37] = -8'd75;
        rom[297][38] = -8'd24;
        rom[297][39] = -8'd20;
        rom[297][40] = -8'd4;
        rom[297][41] = 8'd29;
        rom[297][42] = -8'd36;
        rom[297][43] = 8'd5;
        rom[297][44] = 8'd21;
        rom[297][45] = -8'd19;
        rom[297][46] = 8'd1;
        rom[297][47] = -8'd55;
        rom[297][48] = 8'd1;
        rom[297][49] = -8'd20;
        rom[297][50] = 8'd10;
        rom[297][51] = 8'd15;
        rom[297][52] = 8'd13;
        rom[297][53] = -8'd14;
        rom[297][54] = 8'd0;
        rom[297][55] = -8'd12;
        rom[297][56] = -8'd7;
        rom[297][57] = 8'd38;
        rom[297][58] = -8'd29;
        rom[297][59] = -8'd12;
        rom[297][60] = -8'd20;
        rom[297][61] = -8'd76;
        rom[297][62] = 8'd4;
        rom[297][63] = 8'd8;
        rom[298][0] = 8'd14;
        rom[298][1] = 8'd0;
        rom[298][2] = 8'd18;
        rom[298][3] = -8'd18;
        rom[298][4] = -8'd41;
        rom[298][5] = -8'd14;
        rom[298][6] = -8'd14;
        rom[298][7] = 8'd17;
        rom[298][8] = 8'd5;
        rom[298][9] = 8'd30;
        rom[298][10] = -8'd13;
        rom[298][11] = 8'd19;
        rom[298][12] = 8'd4;
        rom[298][13] = -8'd1;
        rom[298][14] = 8'd16;
        rom[298][15] = -8'd9;
        rom[298][16] = 8'd32;
        rom[298][17] = -8'd35;
        rom[298][18] = 8'd10;
        rom[298][19] = 8'd23;
        rom[298][20] = -8'd5;
        rom[298][21] = 8'd13;
        rom[298][22] = -8'd26;
        rom[298][23] = 8'd0;
        rom[298][24] = -8'd16;
        rom[298][25] = 8'd8;
        rom[298][26] = -8'd5;
        rom[298][27] = 8'd16;
        rom[298][28] = -8'd4;
        rom[298][29] = 8'd0;
        rom[298][30] = 8'd25;
        rom[298][31] = 8'd31;
        rom[298][32] = 8'd13;
        rom[298][33] = 8'd23;
        rom[298][34] = -8'd31;
        rom[298][35] = -8'd26;
        rom[298][36] = -8'd9;
        rom[298][37] = -8'd30;
        rom[298][38] = 8'd4;
        rom[298][39] = 8'd14;
        rom[298][40] = -8'd3;
        rom[298][41] = 8'd12;
        rom[298][42] = 8'd9;
        rom[298][43] = -8'd20;
        rom[298][44] = -8'd18;
        rom[298][45] = -8'd2;
        rom[298][46] = 8'd20;
        rom[298][47] = -8'd28;
        rom[298][48] = 8'd11;
        rom[298][49] = -8'd1;
        rom[298][50] = 8'd21;
        rom[298][51] = -8'd22;
        rom[298][52] = -8'd1;
        rom[298][53] = -8'd38;
        rom[298][54] = -8'd23;
        rom[298][55] = 8'd7;
        rom[298][56] = -8'd18;
        rom[298][57] = 8'd16;
        rom[298][58] = -8'd40;
        rom[298][59] = -8'd5;
        rom[298][60] = -8'd5;
        rom[298][61] = -8'd11;
        rom[298][62] = 8'd13;
        rom[298][63] = 8'd11;
        rom[299][0] = -8'd45;
        rom[299][1] = -8'd40;
        rom[299][2] = -8'd12;
        rom[299][3] = -8'd28;
        rom[299][4] = 8'd10;
        rom[299][5] = -8'd3;
        rom[299][6] = -8'd13;
        rom[299][7] = 8'd3;
        rom[299][8] = 8'd7;
        rom[299][9] = 8'd5;
        rom[299][10] = 8'd44;
        rom[299][11] = -8'd20;
        rom[299][12] = 8'd5;
        rom[299][13] = -8'd16;
        rom[299][14] = -8'd35;
        rom[299][15] = -8'd20;
        rom[299][16] = -8'd19;
        rom[299][17] = -8'd26;
        rom[299][18] = 8'd13;
        rom[299][19] = 8'd4;
        rom[299][20] = -8'd5;
        rom[299][21] = -8'd6;
        rom[299][22] = -8'd61;
        rom[299][23] = -8'd32;
        rom[299][24] = -8'd7;
        rom[299][25] = -8'd52;
        rom[299][26] = -8'd33;
        rom[299][27] = 8'd36;
        rom[299][28] = 8'd13;
        rom[299][29] = -8'd62;
        rom[299][30] = -8'd12;
        rom[299][31] = 8'd2;
        rom[299][32] = -8'd21;
        rom[299][33] = -8'd31;
        rom[299][34] = -8'd24;
        rom[299][35] = -8'd7;
        rom[299][36] = 8'd6;
        rom[299][37] = 8'd6;
        rom[299][38] = 8'd13;
        rom[299][39] = -8'd9;
        rom[299][40] = 8'd9;
        rom[299][41] = 8'd26;
        rom[299][42] = -8'd28;
        rom[299][43] = 8'd26;
        rom[299][44] = -8'd12;
        rom[299][45] = 8'd12;
        rom[299][46] = 8'd16;
        rom[299][47] = 8'd13;
        rom[299][48] = -8'd35;
        rom[299][49] = -8'd24;
        rom[299][50] = -8'd16;
        rom[299][51] = 8'd8;
        rom[299][52] = -8'd34;
        rom[299][53] = 8'd20;
        rom[299][54] = -8'd8;
        rom[299][55] = -8'd8;
        rom[299][56] = -8'd11;
        rom[299][57] = -8'd93;
        rom[299][58] = -8'd19;
        rom[299][59] = 8'd17;
        rom[299][60] = -8'd36;
        rom[299][61] = 8'd10;
        rom[299][62] = -8'd57;
        rom[299][63] = -8'd4;
        rom[300][0] = 8'd6;
        rom[300][1] = -8'd25;
        rom[300][2] = -8'd16;
        rom[300][3] = 8'd5;
        rom[300][4] = -8'd10;
        rom[300][5] = 8'd7;
        rom[300][6] = -8'd3;
        rom[300][7] = 8'd20;
        rom[300][8] = -8'd22;
        rom[300][9] = -8'd50;
        rom[300][10] = -8'd8;
        rom[300][11] = -8'd21;
        rom[300][12] = -8'd13;
        rom[300][13] = 8'd0;
        rom[300][14] = -8'd29;
        rom[300][15] = 8'd10;
        rom[300][16] = -8'd25;
        rom[300][17] = 8'd27;
        rom[300][18] = -8'd3;
        rom[300][19] = -8'd35;
        rom[300][20] = -8'd5;
        rom[300][21] = -8'd15;
        rom[300][22] = -8'd37;
        rom[300][23] = 8'd10;
        rom[300][24] = -8'd4;
        rom[300][25] = -8'd47;
        rom[300][26] = -8'd17;
        rom[300][27] = -8'd2;
        rom[300][28] = -8'd47;
        rom[300][29] = -8'd11;
        rom[300][30] = 8'd16;
        rom[300][31] = -8'd3;
        rom[300][32] = -8'd48;
        rom[300][33] = -8'd23;
        rom[300][34] = -8'd42;
        rom[300][35] = -8'd27;
        rom[300][36] = 8'd24;
        rom[300][37] = 8'd16;
        rom[300][38] = 8'd29;
        rom[300][39] = 8'd36;
        rom[300][40] = -8'd32;
        rom[300][41] = -8'd37;
        rom[300][42] = 8'd11;
        rom[300][43] = 8'd2;
        rom[300][44] = 8'd10;
        rom[300][45] = -8'd24;
        rom[300][46] = 8'd15;
        rom[300][47] = -8'd24;
        rom[300][48] = -8'd19;
        rom[300][49] = 8'd5;
        rom[300][50] = -8'd15;
        rom[300][51] = -8'd25;
        rom[300][52] = -8'd44;
        rom[300][53] = 8'd1;
        rom[300][54] = 8'd12;
        rom[300][55] = 8'd8;
        rom[300][56] = -8'd74;
        rom[300][57] = -8'd12;
        rom[300][58] = -8'd55;
        rom[300][59] = 8'd6;
        rom[300][60] = -8'd19;
        rom[300][61] = -8'd12;
        rom[300][62] = -8'd19;
        rom[300][63] = -8'd6;
        rom[301][0] = 8'd4;
        rom[301][1] = -8'd18;
        rom[301][2] = -8'd20;
        rom[301][3] = 8'd12;
        rom[301][4] = 8'd41;
        rom[301][5] = 8'd9;
        rom[301][6] = 8'd54;
        rom[301][7] = 8'd21;
        rom[301][8] = -8'd55;
        rom[301][9] = 8'd0;
        rom[301][10] = -8'd3;
        rom[301][11] = -8'd18;
        rom[301][12] = -8'd10;
        rom[301][13] = 8'd8;
        rom[301][14] = 8'd3;
        rom[301][15] = -8'd39;
        rom[301][16] = -8'd43;
        rom[301][17] = 8'd1;
        rom[301][18] = -8'd2;
        rom[301][19] = -8'd66;
        rom[301][20] = -8'd7;
        rom[301][21] = -8'd25;
        rom[301][22] = 8'd1;
        rom[301][23] = -8'd63;
        rom[301][24] = 8'd48;
        rom[301][25] = -8'd18;
        rom[301][26] = -8'd42;
        rom[301][27] = 8'd4;
        rom[301][28] = -8'd31;
        rom[301][29] = -8'd32;
        rom[301][30] = 8'd54;
        rom[301][31] = 8'd2;
        rom[301][32] = -8'd65;
        rom[301][33] = -8'd10;
        rom[301][34] = 8'd7;
        rom[301][35] = 8'd4;
        rom[301][36] = 8'd9;
        rom[301][37] = -8'd9;
        rom[301][38] = -8'd17;
        rom[301][39] = -8'd13;
        rom[301][40] = -8'd9;
        rom[301][41] = -8'd39;
        rom[301][42] = 8'd21;
        rom[301][43] = -8'd2;
        rom[301][44] = 8'd8;
        rom[301][45] = -8'd55;
        rom[301][46] = 8'd20;
        rom[301][47] = 8'd16;
        rom[301][48] = 8'd5;
        rom[301][49] = -8'd19;
        rom[301][50] = 8'd8;
        rom[301][51] = -8'd16;
        rom[301][52] = -8'd37;
        rom[301][53] = 8'd14;
        rom[301][54] = -8'd19;
        rom[301][55] = -8'd19;
        rom[301][56] = 8'd6;
        rom[301][57] = -8'd33;
        rom[301][58] = -8'd66;
        rom[301][59] = 8'd36;
        rom[301][60] = 8'd46;
        rom[301][61] = 8'd23;
        rom[301][62] = -8'd29;
        rom[301][63] = -8'd4;
        rom[302][0] = -8'd30;
        rom[302][1] = -8'd29;
        rom[302][2] = -8'd12;
        rom[302][3] = -8'd51;
        rom[302][4] = -8'd16;
        rom[302][5] = -8'd10;
        rom[302][6] = -8'd9;
        rom[302][7] = -8'd32;
        rom[302][8] = -8'd13;
        rom[302][9] = -8'd67;
        rom[302][10] = -8'd40;
        rom[302][11] = -8'd31;
        rom[302][12] = -8'd2;
        rom[302][13] = -8'd7;
        rom[302][14] = -8'd9;
        rom[302][15] = -8'd26;
        rom[302][16] = -8'd43;
        rom[302][17] = -8'd30;
        rom[302][18] = -8'd14;
        rom[302][19] = 8'd23;
        rom[302][20] = -8'd11;
        rom[302][21] = -8'd12;
        rom[302][22] = 8'd2;
        rom[302][23] = -8'd6;
        rom[302][24] = 8'd20;
        rom[302][25] = -8'd39;
        rom[302][26] = 8'd5;
        rom[302][27] = 8'd7;
        rom[302][28] = -8'd20;
        rom[302][29] = 8'd13;
        rom[302][30] = 8'd7;
        rom[302][31] = -8'd23;
        rom[302][32] = 8'd23;
        rom[302][33] = 8'd49;
        rom[302][34] = 8'd17;
        rom[302][35] = 8'd13;
        rom[302][36] = 8'd25;
        rom[302][37] = -8'd6;
        rom[302][38] = -8'd1;
        rom[302][39] = -8'd54;
        rom[302][40] = -8'd11;
        rom[302][41] = 8'd10;
        rom[302][42] = -8'd9;
        rom[302][43] = 8'd11;
        rom[302][44] = -8'd25;
        rom[302][45] = -8'd10;
        rom[302][46] = 8'd11;
        rom[302][47] = -8'd23;
        rom[302][48] = -8'd30;
        rom[302][49] = 8'd26;
        rom[302][50] = -8'd49;
        rom[302][51] = -8'd7;
        rom[302][52] = 8'd13;
        rom[302][53] = -8'd9;
        rom[302][54] = -8'd22;
        rom[302][55] = -8'd10;
        rom[302][56] = 8'd1;
        rom[302][57] = 8'd2;
        rom[302][58] = -8'd10;
        rom[302][59] = -8'd20;
        rom[302][60] = -8'd44;
        rom[302][61] = 8'd1;
        rom[302][62] = -8'd15;
        rom[302][63] = -8'd58;
        rom[303][0] = -8'd24;
        rom[303][1] = 8'd22;
        rom[303][2] = -8'd77;
        rom[303][3] = -8'd9;
        rom[303][4] = -8'd21;
        rom[303][5] = -8'd14;
        rom[303][6] = 8'd3;
        rom[303][7] = -8'd38;
        rom[303][8] = -8'd35;
        rom[303][9] = -8'd65;
        rom[303][10] = 8'd53;
        rom[303][11] = 8'd7;
        rom[303][12] = -8'd1;
        rom[303][13] = -8'd3;
        rom[303][14] = 8'd18;
        rom[303][15] = -8'd57;
        rom[303][16] = -8'd6;
        rom[303][17] = 8'd22;
        rom[303][18] = -8'd35;
        rom[303][19] = 8'd20;
        rom[303][20] = 8'd0;
        rom[303][21] = 8'd26;
        rom[303][22] = 8'd17;
        rom[303][23] = 8'd16;
        rom[303][24] = 8'd27;
        rom[303][25] = -8'd4;
        rom[303][26] = -8'd2;
        rom[303][27] = 8'd17;
        rom[303][28] = -8'd39;
        rom[303][29] = 8'd5;
        rom[303][30] = 8'd8;
        rom[303][31] = 8'd48;
        rom[303][32] = 8'd7;
        rom[303][33] = 8'd25;
        rom[303][34] = 8'd26;
        rom[303][35] = 8'd28;
        rom[303][36] = -8'd24;
        rom[303][37] = 8'd18;
        rom[303][38] = 8'd6;
        rom[303][39] = 8'd35;
        rom[303][40] = 8'd3;
        rom[303][41] = -8'd19;
        rom[303][42] = 8'd10;
        rom[303][43] = -8'd21;
        rom[303][44] = -8'd19;
        rom[303][45] = -8'd14;
        rom[303][46] = -8'd24;
        rom[303][47] = -8'd13;
        rom[303][48] = -8'd3;
        rom[303][49] = 8'd16;
        rom[303][50] = -8'd4;
        rom[303][51] = 8'd11;
        rom[303][52] = -8'd37;
        rom[303][53] = -8'd3;
        rom[303][54] = 8'd29;
        rom[303][55] = 8'd4;
        rom[303][56] = -8'd20;
        rom[303][57] = 8'd31;
        rom[303][58] = -8'd18;
        rom[303][59] = -8'd30;
        rom[303][60] = 8'd5;
        rom[303][61] = 8'd6;
        rom[303][62] = -8'd16;
        rom[303][63] = -8'd17;
        rom[304][0] = -8'd13;
        rom[304][1] = 8'd29;
        rom[304][2] = -8'd58;
        rom[304][3] = -8'd8;
        rom[304][4] = 8'd8;
        rom[304][5] = -8'd47;
        rom[304][6] = 8'd18;
        rom[304][7] = -8'd13;
        rom[304][8] = -8'd18;
        rom[304][9] = -8'd28;
        rom[304][10] = -8'd19;
        rom[304][11] = -8'd12;
        rom[304][12] = 8'd12;
        rom[304][13] = -8'd28;
        rom[304][14] = 8'd14;
        rom[304][15] = 8'd8;
        rom[304][16] = 8'd23;
        rom[304][17] = 8'd41;
        rom[304][18] = 8'd19;
        rom[304][19] = 8'd6;
        rom[304][20] = -8'd1;
        rom[304][21] = 8'd7;
        rom[304][22] = -8'd29;
        rom[304][23] = -8'd29;
        rom[304][24] = 8'd18;
        rom[304][25] = 8'd14;
        rom[304][26] = -8'd44;
        rom[304][27] = -8'd2;
        rom[304][28] = -8'd38;
        rom[304][29] = -8'd53;
        rom[304][30] = 8'd26;
        rom[304][31] = -8'd15;
        rom[304][32] = -8'd2;
        rom[304][33] = 8'd13;
        rom[304][34] = -8'd20;
        rom[304][35] = 8'd2;
        rom[304][36] = 8'd3;
        rom[304][37] = -8'd10;
        rom[304][38] = 8'd5;
        rom[304][39] = -8'd20;
        rom[304][40] = 8'd25;
        rom[304][41] = -8'd13;
        rom[304][42] = -8'd5;
        rom[304][43] = 8'd8;
        rom[304][44] = 8'd3;
        rom[304][45] = 8'd13;
        rom[304][46] = 8'd25;
        rom[304][47] = -8'd4;
        rom[304][48] = 8'd11;
        rom[304][49] = -8'd15;
        rom[304][50] = 8'd16;
        rom[304][51] = -8'd54;
        rom[304][52] = -8'd32;
        rom[304][53] = -8'd11;
        rom[304][54] = 8'd15;
        rom[304][55] = -8'd11;
        rom[304][56] = 8'd15;
        rom[304][57] = -8'd1;
        rom[304][58] = -8'd1;
        rom[304][59] = -8'd6;
        rom[304][60] = -8'd23;
        rom[304][61] = -8'd6;
        rom[304][62] = 8'd23;
        rom[304][63] = -8'd25;
        rom[305][0] = -8'd50;
        rom[305][1] = -8'd31;
        rom[305][2] = -8'd1;
        rom[305][3] = -8'd21;
        rom[305][4] = 8'd10;
        rom[305][5] = 8'd13;
        rom[305][6] = -8'd44;
        rom[305][7] = -8'd25;
        rom[305][8] = 8'd27;
        rom[305][9] = -8'd9;
        rom[305][10] = 8'd14;
        rom[305][11] = 8'd4;
        rom[305][12] = -8'd6;
        rom[305][13] = 8'd66;
        rom[305][14] = -8'd21;
        rom[305][15] = 8'd3;
        rom[305][16] = 8'd10;
        rom[305][17] = 8'd14;
        rom[305][18] = -8'd29;
        rom[305][19] = -8'd12;
        rom[305][20] = 8'd1;
        rom[305][21] = -8'd30;
        rom[305][22] = -8'd21;
        rom[305][23] = 8'd2;
        rom[305][24] = -8'd26;
        rom[305][25] = 8'd10;
        rom[305][26] = -8'd24;
        rom[305][27] = -8'd45;
        rom[305][28] = 8'd27;
        rom[305][29] = -8'd51;
        rom[305][30] = 8'd12;
        rom[305][31] = 8'd3;
        rom[305][32] = -8'd10;
        rom[305][33] = -8'd25;
        rom[305][34] = 8'd7;
        rom[305][35] = -8'd21;
        rom[305][36] = 8'd37;
        rom[305][37] = 8'd7;
        rom[305][38] = -8'd13;
        rom[305][39] = -8'd39;
        rom[305][40] = 8'd1;
        rom[305][41] = 8'd18;
        rom[305][42] = 8'd11;
        rom[305][43] = 8'd20;
        rom[305][44] = 8'd36;
        rom[305][45] = 8'd16;
        rom[305][46] = -8'd3;
        rom[305][47] = 8'd1;
        rom[305][48] = 8'd0;
        rom[305][49] = 8'd22;
        rom[305][50] = -8'd14;
        rom[305][51] = -8'd9;
        rom[305][52] = -8'd22;
        rom[305][53] = 8'd10;
        rom[305][54] = 8'd31;
        rom[305][55] = -8'd16;
        rom[305][56] = 8'd15;
        rom[305][57] = 8'd22;
        rom[305][58] = -8'd13;
        rom[305][59] = 8'd37;
        rom[305][60] = 8'd10;
        rom[305][61] = -8'd17;
        rom[305][62] = -8'd6;
        rom[305][63] = 8'd27;
        rom[306][0] = -8'd4;
        rom[306][1] = 8'd10;
        rom[306][2] = 8'd6;
        rom[306][3] = -8'd36;
        rom[306][4] = -8'd1;
        rom[306][5] = 8'd1;
        rom[306][6] = 8'd8;
        rom[306][7] = -8'd11;
        rom[306][8] = -8'd25;
        rom[306][9] = -8'd18;
        rom[306][10] = 8'd0;
        rom[306][11] = 8'd9;
        rom[306][12] = 8'd5;
        rom[306][13] = 8'd12;
        rom[306][14] = -8'd8;
        rom[306][15] = -8'd29;
        rom[306][16] = -8'd50;
        rom[306][17] = -8'd26;
        rom[306][18] = -8'd33;
        rom[306][19] = 8'd18;
        rom[306][20] = -8'd10;
        rom[306][21] = 8'd10;
        rom[306][22] = 8'd23;
        rom[306][23] = 8'd31;
        rom[306][24] = -8'd30;
        rom[306][25] = -8'd31;
        rom[306][26] = -8'd24;
        rom[306][27] = 8'd8;
        rom[306][28] = -8'd6;
        rom[306][29] = 8'd20;
        rom[306][30] = -8'd11;
        rom[306][31] = -8'd7;
        rom[306][32] = 8'd8;
        rom[306][33] = -8'd12;
        rom[306][34] = 8'd45;
        rom[306][35] = -8'd4;
        rom[306][36] = -8'd9;
        rom[306][37] = 8'd14;
        rom[306][38] = 8'd9;
        rom[306][39] = -8'd30;
        rom[306][40] = -8'd32;
        rom[306][41] = -8'd1;
        rom[306][42] = -8'd33;
        rom[306][43] = 8'd33;
        rom[306][44] = 8'd34;
        rom[306][45] = -8'd61;
        rom[306][46] = -8'd1;
        rom[306][47] = 8'd2;
        rom[306][48] = -8'd9;
        rom[306][49] = -8'd1;
        rom[306][50] = -8'd16;
        rom[306][51] = -8'd11;
        rom[306][52] = 8'd14;
        rom[306][53] = -8'd29;
        rom[306][54] = 8'd12;
        rom[306][55] = -8'd25;
        rom[306][56] = 8'd11;
        rom[306][57] = -8'd18;
        rom[306][58] = 8'd21;
        rom[306][59] = -8'd1;
        rom[306][60] = -8'd25;
        rom[306][61] = 8'd16;
        rom[306][62] = 8'd17;
        rom[306][63] = -8'd14;
        rom[307][0] = 8'd0;
        rom[307][1] = -8'd25;
        rom[307][2] = -8'd19;
        rom[307][3] = -8'd23;
        rom[307][4] = -8'd33;
        rom[307][5] = -8'd28;
        rom[307][6] = -8'd15;
        rom[307][7] = 8'd5;
        rom[307][8] = -8'd1;
        rom[307][9] = -8'd40;
        rom[307][10] = 8'd29;
        rom[307][11] = -8'd9;
        rom[307][12] = -8'd16;
        rom[307][13] = -8'd5;
        rom[307][14] = 8'd9;
        rom[307][15] = -8'd6;
        rom[307][16] = -8'd20;
        rom[307][17] = 8'd13;
        rom[307][18] = -8'd6;
        rom[307][19] = -8'd11;
        rom[307][20] = 8'd0;
        rom[307][21] = 8'd10;
        rom[307][22] = 8'd8;
        rom[307][23] = -8'd26;
        rom[307][24] = 8'd12;
        rom[307][25] = 8'd27;
        rom[307][26] = 8'd8;
        rom[307][27] = -8'd19;
        rom[307][28] = -8'd13;
        rom[307][29] = 8'd14;
        rom[307][30] = -8'd20;
        rom[307][31] = -8'd2;
        rom[307][32] = -8'd5;
        rom[307][33] = -8'd27;
        rom[307][34] = -8'd22;
        rom[307][35] = -8'd17;
        rom[307][36] = -8'd16;
        rom[307][37] = 8'd16;
        rom[307][38] = -8'd11;
        rom[307][39] = 8'd26;
        rom[307][40] = -8'd15;
        rom[307][41] = -8'd34;
        rom[307][42] = -8'd37;
        rom[307][43] = -8'd16;
        rom[307][44] = 8'd3;
        rom[307][45] = -8'd27;
        rom[307][46] = -8'd31;
        rom[307][47] = -8'd26;
        rom[307][48] = 8'd34;
        rom[307][49] = 8'd6;
        rom[307][50] = -8'd35;
        rom[307][51] = -8'd20;
        rom[307][52] = 8'd0;
        rom[307][53] = -8'd20;
        rom[307][54] = -8'd64;
        rom[307][55] = 8'd27;
        rom[307][56] = -8'd32;
        rom[307][57] = -8'd39;
        rom[307][58] = 8'd0;
        rom[307][59] = -8'd4;
        rom[307][60] = 8'd3;
        rom[307][61] = -8'd14;
        rom[307][62] = 8'd35;
        rom[307][63] = -8'd7;
        rom[308][0] = 8'd15;
        rom[308][1] = -8'd43;
        rom[308][2] = -8'd86;
        rom[308][3] = -8'd2;
        rom[308][4] = 8'd30;
        rom[308][5] = -8'd25;
        rom[308][6] = 8'd10;
        rom[308][7] = -8'd18;
        rom[308][8] = -8'd35;
        rom[308][9] = -8'd51;
        rom[308][10] = 8'd15;
        rom[308][11] = -8'd7;
        rom[308][12] = -8'd42;
        rom[308][13] = -8'd49;
        rom[308][14] = -8'd2;
        rom[308][15] = -8'd68;
        rom[308][16] = -8'd32;
        rom[308][17] = 8'd16;
        rom[308][18] = -8'd2;
        rom[308][19] = -8'd30;
        rom[308][20] = -8'd16;
        rom[308][21] = -8'd30;
        rom[308][22] = -8'd35;
        rom[308][23] = 8'd3;
        rom[308][24] = -8'd14;
        rom[308][25] = -8'd11;
        rom[308][26] = -8'd5;
        rom[308][27] = -8'd35;
        rom[308][28] = -8'd21;
        rom[308][29] = -8'd43;
        rom[308][30] = -8'd26;
        rom[308][31] = -8'd8;
        rom[308][32] = -8'd35;
        rom[308][33] = -8'd4;
        rom[308][34] = -8'd24;
        rom[308][35] = 8'd21;
        rom[308][36] = -8'd39;
        rom[308][37] = -8'd15;
        rom[308][38] = -8'd65;
        rom[308][39] = 8'd24;
        rom[308][40] = 8'd3;
        rom[308][41] = 8'd10;
        rom[308][42] = -8'd56;
        rom[308][43] = -8'd91;
        rom[308][44] = 8'd21;
        rom[308][45] = 8'd2;
        rom[308][46] = -8'd11;
        rom[308][47] = -8'd15;
        rom[308][48] = -8'd31;
        rom[308][49] = 8'd14;
        rom[308][50] = -8'd36;
        rom[308][51] = 8'd7;
        rom[308][52] = -8'd26;
        rom[308][53] = 8'd13;
        rom[308][54] = -8'd11;
        rom[308][55] = 8'd11;
        rom[308][56] = 8'd26;
        rom[308][57] = 8'd14;
        rom[308][58] = -8'd23;
        rom[308][59] = -8'd16;
        rom[308][60] = -8'd21;
        rom[308][61] = -8'd11;
        rom[308][62] = -8'd19;
        rom[308][63] = -8'd14;
        rom[309][0] = 8'd9;
        rom[309][1] = -8'd37;
        rom[309][2] = -8'd26;
        rom[309][3] = -8'd65;
        rom[309][4] = -8'd27;
        rom[309][5] = 8'd10;
        rom[309][6] = 8'd18;
        rom[309][7] = 8'd8;
        rom[309][8] = 8'd7;
        rom[309][9] = 8'd13;
        rom[309][10] = -8'd73;
        rom[309][11] = -8'd1;
        rom[309][12] = 8'd18;
        rom[309][13] = 8'd7;
        rom[309][14] = 8'd60;
        rom[309][15] = -8'd8;
        rom[309][16] = 8'd16;
        rom[309][17] = -8'd28;
        rom[309][18] = 8'd35;
        rom[309][19] = -8'd12;
        rom[309][20] = 8'd0;
        rom[309][21] = -8'd27;
        rom[309][22] = 8'd21;
        rom[309][23] = 8'd2;
        rom[309][24] = 8'd18;
        rom[309][25] = 8'd5;
        rom[309][26] = 8'd2;
        rom[309][27] = 8'd7;
        rom[309][28] = 8'd1;
        rom[309][29] = -8'd20;
        rom[309][30] = -8'd33;
        rom[309][31] = -8'd1;
        rom[309][32] = -8'd42;
        rom[309][33] = 8'd9;
        rom[309][34] = -8'd17;
        rom[309][35] = 8'd3;
        rom[309][36] = 8'd2;
        rom[309][37] = 8'd18;
        rom[309][38] = 8'd35;
        rom[309][39] = -8'd5;
        rom[309][40] = 8'd1;
        rom[309][41] = 8'd23;
        rom[309][42] = -8'd15;
        rom[309][43] = -8'd19;
        rom[309][44] = -8'd43;
        rom[309][45] = 8'd0;
        rom[309][46] = 8'd15;
        rom[309][47] = 8'd39;
        rom[309][48] = 8'd8;
        rom[309][49] = -8'd43;
        rom[309][50] = -8'd9;
        rom[309][51] = 8'd7;
        rom[309][52] = -8'd21;
        rom[309][53] = 8'd7;
        rom[309][54] = -8'd6;
        rom[309][55] = -8'd34;
        rom[309][56] = -8'd19;
        rom[309][57] = 8'd0;
        rom[309][58] = 8'd11;
        rom[309][59] = 8'd13;
        rom[309][60] = 8'd29;
        rom[309][61] = 8'd16;
        rom[309][62] = -8'd8;
        rom[309][63] = 8'd16;
        rom[310][0] = 8'd7;
        rom[310][1] = -8'd1;
        rom[310][2] = -8'd1;
        rom[310][3] = 8'd0;
        rom[310][4] = 8'd0;
        rom[310][5] = 8'd7;
        rom[310][6] = -8'd4;
        rom[310][7] = -8'd4;
        rom[310][8] = -8'd3;
        rom[310][9] = 8'd7;
        rom[310][10] = 8'd4;
        rom[310][11] = -8'd4;
        rom[310][12] = 8'd0;
        rom[310][13] = 8'd8;
        rom[310][14] = 8'd9;
        rom[310][15] = -8'd7;
        rom[310][16] = 8'd2;
        rom[310][17] = 8'd3;
        rom[310][18] = 8'd4;
        rom[310][19] = 8'd0;
        rom[310][20] = -8'd2;
        rom[310][21] = -8'd4;
        rom[310][22] = 8'd8;
        rom[310][23] = -8'd3;
        rom[310][24] = 8'd4;
        rom[310][25] = -8'd6;
        rom[310][26] = -8'd12;
        rom[310][27] = -8'd2;
        rom[310][28] = 8'd3;
        rom[310][29] = -8'd9;
        rom[310][30] = 8'd10;
        rom[310][31] = -8'd9;
        rom[310][32] = -8'd10;
        rom[310][33] = -8'd9;
        rom[310][34] = 8'd3;
        rom[310][35] = 8'd5;
        rom[310][36] = -8'd6;
        rom[310][37] = 8'd11;
        rom[310][38] = -8'd11;
        rom[310][39] = 8'd0;
        rom[310][40] = 8'd2;
        rom[310][41] = -8'd8;
        rom[310][42] = -8'd1;
        rom[310][43] = -8'd7;
        rom[310][44] = 8'd5;
        rom[310][45] = -8'd1;
        rom[310][46] = 8'd3;
        rom[310][47] = 8'd6;
        rom[310][48] = 8'd6;
        rom[310][49] = 8'd3;
        rom[310][50] = -8'd4;
        rom[310][51] = 8'd0;
        rom[310][52] = 8'd9;
        rom[310][53] = 8'd5;
        rom[310][54] = -8'd9;
        rom[310][55] = 8'd0;
        rom[310][56] = 8'd1;
        rom[310][57] = -8'd6;
        rom[310][58] = 8'd6;
        rom[310][59] = 8'd6;
        rom[310][60] = 8'd5;
        rom[310][61] = 8'd5;
        rom[310][62] = 8'd6;
        rom[310][63] = 8'd8;
        rom[311][0] = 8'd29;
        rom[311][1] = -8'd50;
        rom[311][2] = -8'd52;
        rom[311][3] = -8'd11;
        rom[311][4] = 8'd45;
        rom[311][5] = -8'd30;
        rom[311][6] = -8'd4;
        rom[311][7] = -8'd1;
        rom[311][8] = -8'd18;
        rom[311][9] = -8'd7;
        rom[311][10] = -8'd18;
        rom[311][11] = -8'd18;
        rom[311][12] = -8'd33;
        rom[311][13] = 8'd12;
        rom[311][14] = 8'd7;
        rom[311][15] = -8'd62;
        rom[311][16] = 8'd4;
        rom[311][17] = 8'd16;
        rom[311][18] = -8'd47;
        rom[311][19] = -8'd56;
        rom[311][20] = -8'd13;
        rom[311][21] = 8'd9;
        rom[311][22] = -8'd36;
        rom[311][23] = 8'd38;
        rom[311][24] = -8'd38;
        rom[311][25] = 8'd19;
        rom[311][26] = -8'd47;
        rom[311][27] = 8'd12;
        rom[311][28] = -8'd37;
        rom[311][29] = 8'd21;
        rom[311][30] = -8'd28;
        rom[311][31] = -8'd2;
        rom[311][32] = -8'd19;
        rom[311][33] = -8'd13;
        rom[311][34] = 8'd11;
        rom[311][35] = -8'd23;
        rom[311][36] = -8'd13;
        rom[311][37] = 8'd20;
        rom[311][38] = -8'd32;
        rom[311][39] = -8'd8;
        rom[311][40] = 8'd30;
        rom[311][41] = -8'd25;
        rom[311][42] = -8'd34;
        rom[311][43] = -8'd11;
        rom[311][44] = 8'd24;
        rom[311][45] = -8'd38;
        rom[311][46] = 8'd9;
        rom[311][47] = -8'd24;
        rom[311][48] = -8'd37;
        rom[311][49] = 8'd28;
        rom[311][50] = 8'd15;
        rom[311][51] = 8'd15;
        rom[311][52] = 8'd0;
        rom[311][53] = -8'd2;
        rom[311][54] = -8'd7;
        rom[311][55] = -8'd75;
        rom[311][56] = -8'd57;
        rom[311][57] = 8'd3;
        rom[311][58] = -8'd1;
        rom[311][59] = -8'd13;
        rom[311][60] = -8'd52;
        rom[311][61] = 8'd10;
        rom[311][62] = 8'd24;
        rom[311][63] = 8'd23;
        rom[312][0] = -8'd8;
        rom[312][1] = -8'd19;
        rom[312][2] = -8'd21;
        rom[312][3] = -8'd50;
        rom[312][4] = -8'd30;
        rom[312][5] = -8'd17;
        rom[312][6] = -8'd13;
        rom[312][7] = -8'd20;
        rom[312][8] = -8'd52;
        rom[312][9] = -8'd9;
        rom[312][10] = 8'd3;
        rom[312][11] = -8'd23;
        rom[312][12] = -8'd33;
        rom[312][13] = -8'd6;
        rom[312][14] = -8'd30;
        rom[312][15] = -8'd21;
        rom[312][16] = 8'd12;
        rom[312][17] = -8'd15;
        rom[312][18] = -8'd20;
        rom[312][19] = -8'd10;
        rom[312][20] = -8'd16;
        rom[312][21] = 8'd12;
        rom[312][22] = -8'd48;
        rom[312][23] = -8'd4;
        rom[312][24] = 8'd12;
        rom[312][25] = -8'd5;
        rom[312][26] = -8'd11;
        rom[312][27] = -8'd45;
        rom[312][28] = -8'd47;
        rom[312][29] = 8'd4;
        rom[312][30] = 8'd4;
        rom[312][31] = -8'd25;
        rom[312][32] = 8'd9;
        rom[312][33] = -8'd50;
        rom[312][34] = -8'd20;
        rom[312][35] = -8'd13;
        rom[312][36] = 8'd6;
        rom[312][37] = 8'd27;
        rom[312][38] = 8'd7;
        rom[312][39] = -8'd3;
        rom[312][40] = -8'd1;
        rom[312][41] = -8'd21;
        rom[312][42] = -8'd27;
        rom[312][43] = -8'd23;
        rom[312][44] = -8'd1;
        rom[312][45] = -8'd68;
        rom[312][46] = 8'd17;
        rom[312][47] = -8'd10;
        rom[312][48] = -8'd20;
        rom[312][49] = -8'd12;
        rom[312][50] = -8'd57;
        rom[312][51] = -8'd31;
        rom[312][52] = 8'd26;
        rom[312][53] = 8'd11;
        rom[312][54] = -8'd23;
        rom[312][55] = 8'd15;
        rom[312][56] = -8'd42;
        rom[312][57] = -8'd12;
        rom[312][58] = -8'd66;
        rom[312][59] = 8'd23;
        rom[312][60] = -8'd9;
        rom[312][61] = 8'd12;
        rom[312][62] = 8'd4;
        rom[312][63] = -8'd25;
        rom[313][0] = 8'd17;
        rom[313][1] = 8'd11;
        rom[313][2] = 8'd48;
        rom[313][3] = 8'd27;
        rom[313][4] = 8'd18;
        rom[313][5] = 8'd5;
        rom[313][6] = 8'd25;
        rom[313][7] = 8'd3;
        rom[313][8] = -8'd5;
        rom[313][9] = 8'd1;
        rom[313][10] = -8'd7;
        rom[313][11] = 8'd2;
        rom[313][12] = 8'd23;
        rom[313][13] = 8'd30;
        rom[313][14] = -8'd19;
        rom[313][15] = 8'd23;
        rom[313][16] = -8'd12;
        rom[313][17] = 8'd16;
        rom[313][18] = 8'd42;
        rom[313][19] = -8'd1;
        rom[313][20] = -8'd7;
        rom[313][21] = -8'd17;
        rom[313][22] = -8'd29;
        rom[313][23] = 8'd13;
        rom[313][24] = 8'd41;
        rom[313][25] = 8'd17;
        rom[313][26] = -8'd3;
        rom[313][27] = 8'd22;
        rom[313][28] = -8'd11;
        rom[313][29] = 8'd11;
        rom[313][30] = 8'd60;
        rom[313][31] = 8'd32;
        rom[313][32] = -8'd29;
        rom[313][33] = -8'd6;
        rom[313][34] = 8'd19;
        rom[313][35] = -8'd20;
        rom[313][36] = -8'd3;
        rom[313][37] = 8'd7;
        rom[313][38] = -8'd23;
        rom[313][39] = 8'd28;
        rom[313][40] = -8'd32;
        rom[313][41] = -8'd22;
        rom[313][42] = 8'd14;
        rom[313][43] = 8'd28;
        rom[313][44] = 8'd16;
        rom[313][45] = -8'd2;
        rom[313][46] = -8'd13;
        rom[313][47] = 8'd27;
        rom[313][48] = -8'd29;
        rom[313][49] = -8'd6;
        rom[313][50] = 8'd1;
        rom[313][51] = -8'd3;
        rom[313][52] = 8'd7;
        rom[313][53] = -8'd41;
        rom[313][54] = -8'd5;
        rom[313][55] = 8'd3;
        rom[313][56] = -8'd5;
        rom[313][57] = -8'd3;
        rom[313][58] = 8'd12;
        rom[313][59] = 8'd1;
        rom[313][60] = 8'd29;
        rom[313][61] = -8'd12;
        rom[313][62] = 8'd8;
        rom[313][63] = 8'd0;
        rom[314][0] = 8'd15;
        rom[314][1] = 8'd22;
        rom[314][2] = 8'd35;
        rom[314][3] = 8'd14;
        rom[314][4] = 8'd1;
        rom[314][5] = -8'd35;
        rom[314][6] = -8'd5;
        rom[314][7] = 8'd4;
        rom[314][8] = -8'd16;
        rom[314][9] = -8'd43;
        rom[314][10] = 8'd42;
        rom[314][11] = -8'd26;
        rom[314][12] = -8'd31;
        rom[314][13] = 8'd4;
        rom[314][14] = -8'd69;
        rom[314][15] = -8'd18;
        rom[314][16] = 8'd15;
        rom[314][17] = 8'd23;
        rom[314][18] = 8'd16;
        rom[314][19] = -8'd35;
        rom[314][20] = -8'd10;
        rom[314][21] = 8'd27;
        rom[314][22] = 8'd35;
        rom[314][23] = 8'd74;
        rom[314][24] = -8'd2;
        rom[314][25] = 8'd20;
        rom[314][26] = -8'd26;
        rom[314][27] = -8'd24;
        rom[314][28] = -8'd26;
        rom[314][29] = -8'd38;
        rom[314][30] = 8'd6;
        rom[314][31] = 8'd12;
        rom[314][32] = -8'd4;
        rom[314][33] = -8'd31;
        rom[314][34] = 8'd9;
        rom[314][35] = -8'd1;
        rom[314][36] = 8'd23;
        rom[314][37] = 8'd43;
        rom[314][38] = -8'd14;
        rom[314][39] = -8'd52;
        rom[314][40] = -8'd23;
        rom[314][41] = -8'd5;
        rom[314][42] = -8'd11;
        rom[314][43] = -8'd17;
        rom[314][44] = -8'd4;
        rom[314][45] = -8'd69;
        rom[314][46] = 8'd14;
        rom[314][47] = -8'd17;
        rom[314][48] = 8'd20;
        rom[314][49] = 8'd24;
        rom[314][50] = -8'd67;
        rom[314][51] = 8'd7;
        rom[314][52] = -8'd30;
        rom[314][53] = 8'd14;
        rom[314][54] = 8'd15;
        rom[314][55] = -8'd16;
        rom[314][56] = 8'd38;
        rom[314][57] = -8'd34;
        rom[314][58] = 8'd33;
        rom[314][59] = -8'd24;
        rom[314][60] = 8'd1;
        rom[314][61] = 8'd20;
        rom[314][62] = 8'd8;
        rom[314][63] = -8'd18;
        rom[315][0] = -8'd30;
        rom[315][1] = 8'd10;
        rom[315][2] = -8'd30;
        rom[315][3] = -8'd15;
        rom[315][4] = -8'd16;
        rom[315][5] = -8'd30;
        rom[315][6] = -8'd33;
        rom[315][7] = -8'd3;
        rom[315][8] = -8'd12;
        rom[315][9] = -8'd12;
        rom[315][10] = 8'd31;
        rom[315][11] = -8'd16;
        rom[315][12] = 8'd9;
        rom[315][13] = 8'd12;
        rom[315][14] = 8'd9;
        rom[315][15] = -8'd35;
        rom[315][16] = 8'd44;
        rom[315][17] = 8'd19;
        rom[315][18] = 8'd6;
        rom[315][19] = -8'd3;
        rom[315][20] = -8'd4;
        rom[315][21] = -8'd10;
        rom[315][22] = -8'd17;
        rom[315][23] = -8'd3;
        rom[315][24] = -8'd14;
        rom[315][25] = -8'd55;
        rom[315][26] = 8'd2;
        rom[315][27] = 8'd6;
        rom[315][28] = -8'd19;
        rom[315][29] = -8'd20;
        rom[315][30] = -8'd1;
        rom[315][31] = -8'd31;
        rom[315][32] = -8'd3;
        rom[315][33] = -8'd9;
        rom[315][34] = 8'd19;
        rom[315][35] = -8'd11;
        rom[315][36] = -8'd10;
        rom[315][37] = 8'd8;
        rom[315][38] = -8'd14;
        rom[315][39] = -8'd24;
        rom[315][40] = 8'd5;
        rom[315][41] = -8'd30;
        rom[315][42] = -8'd29;
        rom[315][43] = -8'd22;
        rom[315][44] = 8'd1;
        rom[315][45] = 8'd13;
        rom[315][46] = -8'd18;
        rom[315][47] = 8'd36;
        rom[315][48] = 8'd24;
        rom[315][49] = 8'd12;
        rom[315][50] = -8'd62;
        rom[315][51] = 8'd9;
        rom[315][52] = -8'd39;
        rom[315][53] = -8'd6;
        rom[315][54] = -8'd8;
        rom[315][55] = -8'd38;
        rom[315][56] = -8'd27;
        rom[315][57] = -8'd60;
        rom[315][58] = 8'd15;
        rom[315][59] = -8'd21;
        rom[315][60] = -8'd4;
        rom[315][61] = -8'd22;
        rom[315][62] = -8'd45;
        rom[315][63] = -8'd5;
        rom[316][0] = 8'd0;
        rom[316][1] = 8'd25;
        rom[316][2] = 8'd2;
        rom[316][3] = 8'd0;
        rom[316][4] = 8'd3;
        rom[316][5] = -8'd13;
        rom[316][6] = -8'd15;
        rom[316][7] = 8'd8;
        rom[316][8] = 8'd17;
        rom[316][9] = -8'd19;
        rom[316][10] = -8'd45;
        rom[316][11] = 8'd13;
        rom[316][12] = 8'd19;
        rom[316][13] = -8'd72;
        rom[316][14] = -8'd20;
        rom[316][15] = 8'd21;
        rom[316][16] = 8'd22;
        rom[316][17] = 8'd12;
        rom[316][18] = 8'd13;
        rom[316][19] = -8'd32;
        rom[316][20] = -8'd12;
        rom[316][21] = -8'd52;
        rom[316][22] = -8'd12;
        rom[316][23] = 8'd7;
        rom[316][24] = 8'd3;
        rom[316][25] = 8'd42;
        rom[316][26] = 8'd42;
        rom[316][27] = -8'd32;
        rom[316][28] = -8'd9;
        rom[316][29] = 8'd44;
        rom[316][30] = -8'd10;
        rom[316][31] = 8'd16;
        rom[316][32] = 8'd13;
        rom[316][33] = -8'd24;
        rom[316][34] = -8'd23;
        rom[316][35] = -8'd17;
        rom[316][36] = 8'd4;
        rom[316][37] = 8'd21;
        rom[316][38] = 8'd8;
        rom[316][39] = 8'd12;
        rom[316][40] = -8'd8;
        rom[316][41] = 8'd3;
        rom[316][42] = -8'd35;
        rom[316][43] = 8'd9;
        rom[316][44] = 8'd5;
        rom[316][45] = 8'd27;
        rom[316][46] = -8'd6;
        rom[316][47] = -8'd36;
        rom[316][48] = -8'd4;
        rom[316][49] = -8'd17;
        rom[316][50] = -8'd7;
        rom[316][51] = -8'd14;
        rom[316][52] = -8'd64;
        rom[316][53] = -8'd48;
        rom[316][54] = -8'd25;
        rom[316][55] = 8'd25;
        rom[316][56] = 8'd4;
        rom[316][57] = -8'd21;
        rom[316][58] = -8'd6;
        rom[316][59] = -8'd14;
        rom[316][60] = -8'd21;
        rom[316][61] = -8'd18;
        rom[316][62] = 8'd19;
        rom[316][63] = 8'd14;
        rom[317][0] = 8'd19;
        rom[317][1] = 8'd7;
        rom[317][2] = -8'd4;
        rom[317][3] = -8'd24;
        rom[317][4] = -8'd3;
        rom[317][5] = 8'd4;
        rom[317][6] = -8'd14;
        rom[317][7] = 8'd7;
        rom[317][8] = -8'd5;
        rom[317][9] = 8'd14;
        rom[317][10] = 8'd17;
        rom[317][11] = 8'd3;
        rom[317][12] = -8'd34;
        rom[317][13] = 8'd11;
        rom[317][14] = -8'd37;
        rom[317][15] = 8'd4;
        rom[317][16] = 8'd15;
        rom[317][17] = -8'd39;
        rom[317][18] = 8'd42;
        rom[317][19] = -8'd8;
        rom[317][20] = 8'd3;
        rom[317][21] = 8'd27;
        rom[317][22] = 8'd2;
        rom[317][23] = -8'd18;
        rom[317][24] = 8'd39;
        rom[317][25] = -8'd38;
        rom[317][26] = 8'd4;
        rom[317][27] = -8'd21;
        rom[317][28] = -8'd23;
        rom[317][29] = 8'd19;
        rom[317][30] = -8'd2;
        rom[317][31] = -8'd33;
        rom[317][32] = 8'd14;
        rom[317][33] = 8'd11;
        rom[317][34] = 8'd13;
        rom[317][35] = 8'd0;
        rom[317][36] = 8'd0;
        rom[317][37] = 8'd14;
        rom[317][38] = -8'd25;
        rom[317][39] = -8'd14;
        rom[317][40] = -8'd10;
        rom[317][41] = 8'd16;
        rom[317][42] = 8'd13;
        rom[317][43] = 8'd12;
        rom[317][44] = 8'd29;
        rom[317][45] = -8'd25;
        rom[317][46] = 8'd26;
        rom[317][47] = 8'd35;
        rom[317][48] = 8'd7;
        rom[317][49] = 8'd40;
        rom[317][50] = 8'd21;
        rom[317][51] = -8'd13;
        rom[317][52] = 8'd11;
        rom[317][53] = -8'd13;
        rom[317][54] = 8'd15;
        rom[317][55] = 8'd11;
        rom[317][56] = -8'd44;
        rom[317][57] = -8'd12;
        rom[317][58] = -8'd13;
        rom[317][59] = 8'd33;
        rom[317][60] = -8'd1;
        rom[317][61] = -8'd30;
        rom[317][62] = -8'd22;
        rom[317][63] = 8'd4;
        rom[318][0] = 8'd16;
        rom[318][1] = -8'd29;
        rom[318][2] = -8'd51;
        rom[318][3] = 8'd20;
        rom[318][4] = -8'd17;
        rom[318][5] = 8'd10;
        rom[318][6] = -8'd40;
        rom[318][7] = -8'd7;
        rom[318][8] = -8'd16;
        rom[318][9] = -8'd14;
        rom[318][10] = 8'd13;
        rom[318][11] = 8'd8;
        rom[318][12] = -8'd19;
        rom[318][13] = 8'd2;
        rom[318][14] = -8'd17;
        rom[318][15] = 8'd14;
        rom[318][16] = 8'd23;
        rom[318][17] = 8'd65;
        rom[318][18] = 8'd11;
        rom[318][19] = -8'd9;
        rom[318][20] = -8'd1;
        rom[318][21] = 8'd17;
        rom[318][22] = -8'd61;
        rom[318][23] = -8'd20;
        rom[318][24] = -8'd31;
        rom[318][25] = 8'd37;
        rom[318][26] = -8'd19;
        rom[318][27] = -8'd9;
        rom[318][28] = 8'd2;
        rom[318][29] = -8'd35;
        rom[318][30] = -8'd17;
        rom[318][31] = -8'd13;
        rom[318][32] = -8'd30;
        rom[318][33] = -8'd1;
        rom[318][34] = 8'd16;
        rom[318][35] = 8'd9;
        rom[318][36] = 8'd10;
        rom[318][37] = -8'd3;
        rom[318][38] = -8'd6;
        rom[318][39] = -8'd1;
        rom[318][40] = -8'd14;
        rom[318][41] = -8'd29;
        rom[318][42] = -8'd4;
        rom[318][43] = -8'd46;
        rom[318][44] = 8'd11;
        rom[318][45] = -8'd8;
        rom[318][46] = -8'd6;
        rom[318][47] = 8'd44;
        rom[318][48] = -8'd26;
        rom[318][49] = -8'd38;
        rom[318][50] = 8'd2;
        rom[318][51] = 8'd11;
        rom[318][52] = -8'd25;
        rom[318][53] = 8'd31;
        rom[318][54] = -8'd42;
        rom[318][55] = 8'd32;
        rom[318][56] = -8'd6;
        rom[318][57] = 8'd16;
        rom[318][58] = -8'd25;
        rom[318][59] = -8'd4;
        rom[318][60] = -8'd6;
        rom[318][61] = -8'd11;
        rom[318][62] = 8'd4;
        rom[318][63] = 8'd11;
        rom[319][0] = -8'd11;
        rom[319][1] = -8'd2;
        rom[319][2] = 8'd1;
        rom[319][3] = -8'd29;
        rom[319][4] = -8'd39;
        rom[319][5] = 8'd24;
        rom[319][6] = 8'd5;
        rom[319][7] = -8'd34;
        rom[319][8] = -8'd32;
        rom[319][9] = -8'd46;
        rom[319][10] = -8'd22;
        rom[319][11] = 8'd41;
        rom[319][12] = -8'd6;
        rom[319][13] = -8'd16;
        rom[319][14] = -8'd22;
        rom[319][15] = 8'd18;
        rom[319][16] = -8'd48;
        rom[319][17] = 8'd19;
        rom[319][18] = -8'd5;
        rom[319][19] = -8'd11;
        rom[319][20] = -8'd6;
        rom[319][21] = -8'd13;
        rom[319][22] = 8'd0;
        rom[319][23] = 8'd37;
        rom[319][24] = -8'd14;
        rom[319][25] = 8'd11;
        rom[319][26] = 8'd12;
        rom[319][27] = 8'd3;
        rom[319][28] = 8'd3;
        rom[319][29] = 8'd5;
        rom[319][30] = -8'd47;
        rom[319][31] = -8'd16;
        rom[319][32] = 8'd38;
        rom[319][33] = 8'd21;
        rom[319][34] = 8'd7;
        rom[319][35] = -8'd16;
        rom[319][36] = -8'd17;
        rom[319][37] = 8'd32;
        rom[319][38] = 8'd12;
        rom[319][39] = 8'd23;
        rom[319][40] = 8'd4;
        rom[319][41] = 8'd9;
        rom[319][42] = -8'd17;
        rom[319][43] = -8'd41;
        rom[319][44] = 8'd17;
        rom[319][45] = -8'd19;
        rom[319][46] = -8'd3;
        rom[319][47] = 8'd16;
        rom[319][48] = 8'd17;
        rom[319][49] = -8'd32;
        rom[319][50] = -8'd24;
        rom[319][51] = 8'd3;
        rom[319][52] = -8'd10;
        rom[319][53] = 8'd17;
        rom[319][54] = -8'd34;
        rom[319][55] = -8'd6;
        rom[319][56] = 8'd25;
        rom[319][57] = -8'd29;
        rom[319][58] = 8'd16;
        rom[319][59] = -8'd67;
        rom[319][60] = 8'd7;
        rom[319][61] = -8'd7;
        rom[319][62] = -8'd35;
        rom[319][63] = -8'd14;
        rom[320][0] = -8'd36;
        rom[320][1] = 8'd6;
        rom[320][2] = -8'd14;
        rom[320][3] = -8'd45;
        rom[320][4] = -8'd44;
        rom[320][5] = -8'd65;
        rom[320][6] = 8'd38;
        rom[320][7] = 8'd11;
        rom[320][8] = 8'd11;
        rom[320][9] = 8'd3;
        rom[320][10] = -8'd27;
        rom[320][11] = 8'd6;
        rom[320][12] = 8'd1;
        rom[320][13] = -8'd1;
        rom[320][14] = -8'd14;
        rom[320][15] = 8'd9;
        rom[320][16] = -8'd8;
        rom[320][17] = 8'd10;
        rom[320][18] = 8'd23;
        rom[320][19] = -8'd12;
        rom[320][20] = -8'd16;
        rom[320][21] = 8'd14;
        rom[320][22] = 8'd15;
        rom[320][23] = -8'd36;
        rom[320][24] = -8'd42;
        rom[320][25] = 8'd5;
        rom[320][26] = -8'd38;
        rom[320][27] = -8'd31;
        rom[320][28] = -8'd8;
        rom[320][29] = 8'd13;
        rom[320][30] = -8'd13;
        rom[320][31] = -8'd10;
        rom[320][32] = -8'd34;
        rom[320][33] = -8'd1;
        rom[320][34] = 8'd19;
        rom[320][35] = -8'd13;
        rom[320][36] = -8'd16;
        rom[320][37] = 8'd11;
        rom[320][38] = 8'd7;
        rom[320][39] = 8'd18;
        rom[320][40] = -8'd5;
        rom[320][41] = -8'd20;
        rom[320][42] = -8'd25;
        rom[320][43] = 8'd5;
        rom[320][44] = 8'd12;
        rom[320][45] = 8'd27;
        rom[320][46] = 8'd1;
        rom[320][47] = 8'd31;
        rom[320][48] = -8'd7;
        rom[320][49] = 8'd28;
        rom[320][50] = 8'd14;
        rom[320][51] = -8'd24;
        rom[320][52] = 8'd2;
        rom[320][53] = 8'd16;
        rom[320][54] = -8'd16;
        rom[320][55] = 8'd27;
        rom[320][56] = -8'd11;
        rom[320][57] = 8'd24;
        rom[320][58] = -8'd19;
        rom[320][59] = 8'd0;
        rom[320][60] = 8'd17;
        rom[320][61] = 8'd36;
        rom[320][62] = 8'd12;
        rom[320][63] = -8'd1;
        rom[321][0] = -8'd10;
        rom[321][1] = 8'd15;
        rom[321][2] = -8'd15;
        rom[321][3] = 8'd17;
        rom[321][4] = -8'd28;
        rom[321][5] = 8'd23;
        rom[321][6] = 8'd25;
        rom[321][7] = -8'd3;
        rom[321][8] = 8'd6;
        rom[321][9] = -8'd23;
        rom[321][10] = -8'd35;
        rom[321][11] = 8'd17;
        rom[321][12] = 8'd8;
        rom[321][13] = -8'd89;
        rom[321][14] = 8'd9;
        rom[321][15] = 8'd5;
        rom[321][16] = 8'd17;
        rom[321][17] = 8'd20;
        rom[321][18] = 8'd14;
        rom[321][19] = -8'd77;
        rom[321][20] = -8'd6;
        rom[321][21] = 8'd8;
        rom[321][22] = -8'd64;
        rom[321][23] = -8'd12;
        rom[321][24] = 8'd17;
        rom[321][25] = 8'd1;
        rom[321][26] = 8'd9;
        rom[321][27] = -8'd43;
        rom[321][28] = -8'd23;
        rom[321][29] = 8'd10;
        rom[321][30] = 8'd14;
        rom[321][31] = -8'd11;
        rom[321][32] = 8'd13;
        rom[321][33] = 8'd13;
        rom[321][34] = -8'd9;
        rom[321][35] = -8'd25;
        rom[321][36] = -8'd27;
        rom[321][37] = -8'd29;
        rom[321][38] = 8'd22;
        rom[321][39] = -8'd18;
        rom[321][40] = -8'd21;
        rom[321][41] = -8'd2;
        rom[321][42] = -8'd5;
        rom[321][43] = 8'd7;
        rom[321][44] = -8'd3;
        rom[321][45] = 8'd41;
        rom[321][46] = 8'd4;
        rom[321][47] = -8'd53;
        rom[321][48] = -8'd65;
        rom[321][49] = -8'd4;
        rom[321][50] = -8'd25;
        rom[321][51] = -8'd12;
        rom[321][52] = 8'd3;
        rom[321][53] = -8'd43;
        rom[321][54] = 8'd7;
        rom[321][55] = -8'd30;
        rom[321][56] = -8'd55;
        rom[321][57] = 8'd24;
        rom[321][58] = 8'd28;
        rom[321][59] = 8'd27;
        rom[321][60] = 8'd7;
        rom[321][61] = -8'd7;
        rom[321][62] = -8'd4;
        rom[321][63] = 8'd18;
        rom[322][0] = -8'd22;
        rom[322][1] = -8'd48;
        rom[322][2] = -8'd33;
        rom[322][3] = 8'd11;
        rom[322][4] = -8'd16;
        rom[322][5] = 8'd22;
        rom[322][6] = -8'd58;
        rom[322][7] = -8'd34;
        rom[322][8] = 8'd9;
        rom[322][9] = 8'd20;
        rom[322][10] = 8'd9;
        rom[322][11] = 8'd8;
        rom[322][12] = -8'd41;
        rom[322][13] = 8'd15;
        rom[322][14] = 8'd8;
        rom[322][15] = -8'd62;
        rom[322][16] = -8'd15;
        rom[322][17] = 8'd23;
        rom[322][18] = -8'd14;
        rom[322][19] = -8'd21;
        rom[322][20] = 8'd10;
        rom[322][21] = 8'd28;
        rom[322][22] = -8'd17;
        rom[322][23] = -8'd47;
        rom[322][24] = 8'd17;
        rom[322][25] = -8'd62;
        rom[322][26] = -8'd8;
        rom[322][27] = -8'd33;
        rom[322][28] = -8'd6;
        rom[322][29] = 8'd7;
        rom[322][30] = 8'd10;
        rom[322][31] = -8'd13;
        rom[322][32] = -8'd113;
        rom[322][33] = -8'd57;
        rom[322][34] = -8'd21;
        rom[322][35] = -8'd71;
        rom[322][36] = -8'd6;
        rom[322][37] = -8'd2;
        rom[322][38] = 8'd6;
        rom[322][39] = 8'd4;
        rom[322][40] = 8'd23;
        rom[322][41] = -8'd34;
        rom[322][42] = -8'd59;
        rom[322][43] = -8'd14;
        rom[322][44] = 8'd18;
        rom[322][45] = -8'd4;
        rom[322][46] = -8'd16;
        rom[322][47] = -8'd6;
        rom[322][48] = 8'd6;
        rom[322][49] = -8'd25;
        rom[322][50] = 8'd10;
        rom[322][51] = -8'd24;
        rom[322][52] = 8'd41;
        rom[322][53] = -8'd26;
        rom[322][54] = -8'd78;
        rom[322][55] = -8'd3;
        rom[322][56] = -8'd52;
        rom[322][57] = 8'd5;
        rom[322][58] = -8'd18;
        rom[322][59] = 8'd3;
        rom[322][60] = -8'd58;
        rom[322][61] = 8'd18;
        rom[322][62] = 8'd19;
        rom[322][63] = -8'd47;
        rom[323][0] = -8'd20;
        rom[323][1] = 8'd5;
        rom[323][2] = -8'd9;
        rom[323][3] = -8'd18;
        rom[323][4] = -8'd20;
        rom[323][5] = -8'd22;
        rom[323][6] = 8'd32;
        rom[323][7] = 8'd16;
        rom[323][8] = 8'd3;
        rom[323][9] = 8'd18;
        rom[323][10] = -8'd65;
        rom[323][11] = -8'd36;
        rom[323][12] = 8'd25;
        rom[323][13] = -8'd8;
        rom[323][14] = 8'd3;
        rom[323][15] = 8'd17;
        rom[323][16] = -8'd50;
        rom[323][17] = -8'd32;
        rom[323][18] = 8'd14;
        rom[323][19] = 8'd21;
        rom[323][20] = -8'd8;
        rom[323][21] = 8'd15;
        rom[323][22] = 8'd27;
        rom[323][23] = 8'd4;
        rom[323][24] = -8'd8;
        rom[323][25] = 8'd17;
        rom[323][26] = -8'd43;
        rom[323][27] = -8'd23;
        rom[323][28] = -8'd12;
        rom[323][29] = 8'd15;
        rom[323][30] = 8'd33;
        rom[323][31] = -8'd35;
        rom[323][32] = 8'd12;
        rom[323][33] = -8'd10;
        rom[323][34] = -8'd43;
        rom[323][35] = 8'd32;
        rom[323][36] = 8'd11;
        rom[323][37] = -8'd47;
        rom[323][38] = 8'd21;
        rom[323][39] = 8'd30;
        rom[323][40] = 8'd1;
        rom[323][41] = -8'd2;
        rom[323][42] = 8'd6;
        rom[323][43] = 8'd12;
        rom[323][44] = -8'd36;
        rom[323][45] = -8'd29;
        rom[323][46] = 8'd5;
        rom[323][47] = -8'd52;
        rom[323][48] = -8'd31;
        rom[323][49] = 8'd8;
        rom[323][50] = -8'd30;
        rom[323][51] = 8'd20;
        rom[323][52] = 8'd34;
        rom[323][53] = -8'd15;
        rom[323][54] = -8'd28;
        rom[323][55] = 8'd18;
        rom[323][56] = 8'd7;
        rom[323][57] = -8'd62;
        rom[323][58] = -8'd10;
        rom[323][59] = -8'd9;
        rom[323][60] = 8'd36;
        rom[323][61] = 8'd0;
        rom[323][62] = 8'd5;
        rom[323][63] = 8'd21;
        rom[324][0] = -8'd45;
        rom[324][1] = -8'd10;
        rom[324][2] = -8'd9;
        rom[324][3] = 8'd4;
        rom[324][4] = 8'd9;
        rom[324][5] = -8'd19;
        rom[324][6] = -8'd22;
        rom[324][7] = -8'd63;
        rom[324][8] = 8'd20;
        rom[324][9] = -8'd3;
        rom[324][10] = -8'd53;
        rom[324][11] = -8'd63;
        rom[324][12] = -8'd7;
        rom[324][13] = -8'd10;
        rom[324][14] = 8'd5;
        rom[324][15] = 8'd9;
        rom[324][16] = -8'd14;
        rom[324][17] = 8'd5;
        rom[324][18] = 8'd36;
        rom[324][19] = 8'd12;
        rom[324][20] = -8'd10;
        rom[324][21] = -8'd18;
        rom[324][22] = -8'd20;
        rom[324][23] = 8'd20;
        rom[324][24] = -8'd52;
        rom[324][25] = -8'd12;
        rom[324][26] = -8'd8;
        rom[324][27] = -8'd40;
        rom[324][28] = -8'd25;
        rom[324][29] = 8'd0;
        rom[324][30] = 8'd30;
        rom[324][31] = 8'd4;
        rom[324][32] = 8'd6;
        rom[324][33] = 8'd33;
        rom[324][34] = -8'd50;
        rom[324][35] = -8'd13;
        rom[324][36] = -8'd16;
        rom[324][37] = 8'd26;
        rom[324][38] = -8'd108;
        rom[324][39] = 8'd7;
        rom[324][40] = -8'd21;
        rom[324][41] = -8'd16;
        rom[324][42] = 8'd23;
        rom[324][43] = -8'd4;
        rom[324][44] = -8'd5;
        rom[324][45] = -8'd30;
        rom[324][46] = -8'd3;
        rom[324][47] = 8'd16;
        rom[324][48] = -8'd10;
        rom[324][49] = -8'd10;
        rom[324][50] = -8'd14;
        rom[324][51] = -8'd5;
        rom[324][52] = -8'd15;
        rom[324][53] = 8'd7;
        rom[324][54] = -8'd5;
        rom[324][55] = -8'd2;
        rom[324][56] = 8'd27;
        rom[324][57] = 8'd1;
        rom[324][58] = 8'd25;
        rom[324][59] = -8'd19;
        rom[324][60] = -8'd12;
        rom[324][61] = 8'd8;
        rom[324][62] = -8'd9;
        rom[324][63] = -8'd28;
        rom[325][0] = 8'd1;
        rom[325][1] = -8'd5;
        rom[325][2] = 8'd5;
        rom[325][3] = 8'd3;
        rom[325][4] = 8'd9;
        rom[325][5] = 8'd6;
        rom[325][6] = -8'd8;
        rom[325][7] = 8'd4;
        rom[325][8] = 8'd5;
        rom[325][9] = 8'd9;
        rom[325][10] = 8'd3;
        rom[325][11] = -8'd2;
        rom[325][12] = -8'd4;
        rom[325][13] = -8'd8;
        rom[325][14] = -8'd3;
        rom[325][15] = 8'd12;
        rom[325][16] = 8'd8;
        rom[325][17] = -8'd7;
        rom[325][18] = 8'd6;
        rom[325][19] = -8'd3;
        rom[325][20] = -8'd4;
        rom[325][21] = -8'd4;
        rom[325][22] = 8'd9;
        rom[325][23] = 8'd8;
        rom[325][24] = -8'd9;
        rom[325][25] = -8'd3;
        rom[325][26] = 8'd0;
        rom[325][27] = 8'd7;
        rom[325][28] = 8'd12;
        rom[325][29] = 8'd6;
        rom[325][30] = 8'd8;
        rom[325][31] = -8'd2;
        rom[325][32] = -8'd5;
        rom[325][33] = 8'd1;
        rom[325][34] = -8'd6;
        rom[325][35] = 8'd0;
        rom[325][36] = 8'd8;
        rom[325][37] = -8'd6;
        rom[325][38] = 8'd5;
        rom[325][39] = 8'd0;
        rom[325][40] = 8'd8;
        rom[325][41] = 8'd9;
        rom[325][42] = -8'd8;
        rom[325][43] = 8'd0;
        rom[325][44] = -8'd3;
        rom[325][45] = 8'd4;
        rom[325][46] = -8'd3;
        rom[325][47] = -8'd3;
        rom[325][48] = 8'd4;
        rom[325][49] = 8'd4;
        rom[325][50] = -8'd3;
        rom[325][51] = -8'd6;
        rom[325][52] = 8'd4;
        rom[325][53] = 8'd0;
        rom[325][54] = 8'd0;
        rom[325][55] = -8'd2;
        rom[325][56] = 8'd3;
        rom[325][57] = -8'd6;
        rom[325][58] = -8'd1;
        rom[325][59] = 8'd1;
        rom[325][60] = 8'd0;
        rom[325][61] = 8'd4;
        rom[325][62] = 8'd7;
        rom[325][63] = -8'd6;
        rom[326][0] = -8'd7;
        rom[326][1] = -8'd70;
        rom[326][2] = 8'd7;
        rom[326][3] = 8'd12;
        rom[326][4] = 8'd6;
        rom[326][5] = -8'd42;
        rom[326][6] = -8'd39;
        rom[326][7] = -8'd13;
        rom[326][8] = -8'd6;
        rom[326][9] = 8'd17;
        rom[326][10] = -8'd37;
        rom[326][11] = 8'd20;
        rom[326][12] = -8'd47;
        rom[326][13] = -8'd19;
        rom[326][14] = -8'd8;
        rom[326][15] = -8'd16;
        rom[326][16] = -8'd7;
        rom[326][17] = 8'd19;
        rom[326][18] = -8'd15;
        rom[326][19] = 8'd14;
        rom[326][20] = -8'd12;
        rom[326][21] = 8'd4;
        rom[326][22] = 8'd15;
        rom[326][23] = -8'd9;
        rom[326][24] = -8'd8;
        rom[326][25] = -8'd2;
        rom[326][26] = -8'd33;
        rom[326][27] = -8'd45;
        rom[326][28] = 8'd24;
        rom[326][29] = -8'd19;
        rom[326][30] = 8'd10;
        rom[326][31] = -8'd21;
        rom[326][32] = 8'd14;
        rom[326][33] = 8'd14;
        rom[326][34] = -8'd2;
        rom[326][35] = -8'd27;
        rom[326][36] = -8'd30;
        rom[326][37] = 8'd5;
        rom[326][38] = 8'd7;
        rom[326][39] = -8'd16;
        rom[326][40] = -8'd25;
        rom[326][41] = -8'd11;
        rom[326][42] = 8'd15;
        rom[326][43] = 8'd3;
        rom[326][44] = -8'd10;
        rom[326][45] = -8'd31;
        rom[326][46] = -8'd52;
        rom[326][47] = -8'd32;
        rom[326][48] = 8'd30;
        rom[326][49] = 8'd2;
        rom[326][50] = -8'd3;
        rom[326][51] = -8'd5;
        rom[326][52] = -8'd16;
        rom[326][53] = 8'd39;
        rom[326][54] = 8'd16;
        rom[326][55] = -8'd74;
        rom[326][56] = -8'd18;
        rom[326][57] = 8'd24;
        rom[326][58] = -8'd18;
        rom[326][59] = -8'd19;
        rom[326][60] = 8'd10;
        rom[326][61] = -8'd2;
        rom[326][62] = -8'd18;
        rom[326][63] = 8'd11;
        rom[327][0] = 8'd32;
        rom[327][1] = -8'd22;
        rom[327][2] = -8'd32;
        rom[327][3] = 8'd5;
        rom[327][4] = 8'd7;
        rom[327][5] = -8'd22;
        rom[327][6] = -8'd10;
        rom[327][7] = -8'd32;
        rom[327][8] = 8'd11;
        rom[327][9] = -8'd58;
        rom[327][10] = -8'd21;
        rom[327][11] = -8'd13;
        rom[327][12] = 8'd6;
        rom[327][13] = 8'd16;
        rom[327][14] = -8'd16;
        rom[327][15] = -8'd1;
        rom[327][16] = 8'd6;
        rom[327][17] = 8'd24;
        rom[327][18] = -8'd1;
        rom[327][19] = -8'd45;
        rom[327][20] = 8'd12;
        rom[327][21] = -8'd28;
        rom[327][22] = 8'd60;
        rom[327][23] = 8'd29;
        rom[327][24] = -8'd4;
        rom[327][25] = -8'd24;
        rom[327][26] = 8'd37;
        rom[327][27] = 8'd30;
        rom[327][28] = -8'd6;
        rom[327][29] = 8'd7;
        rom[327][30] = -8'd14;
        rom[327][31] = 8'd14;
        rom[327][32] = -8'd21;
        rom[327][33] = 8'd10;
        rom[327][34] = -8'd15;
        rom[327][35] = -8'd2;
        rom[327][36] = 8'd18;
        rom[327][37] = -8'd21;
        rom[327][38] = 8'd12;
        rom[327][39] = -8'd25;
        rom[327][40] = 8'd3;
        rom[327][41] = 8'd9;
        rom[327][42] = 8'd33;
        rom[327][43] = 8'd11;
        rom[327][44] = -8'd7;
        rom[327][45] = -8'd27;
        rom[327][46] = -8'd7;
        rom[327][47] = 8'd1;
        rom[327][48] = -8'd1;
        rom[327][49] = -8'd38;
        rom[327][50] = 8'd11;
        rom[327][51] = -8'd43;
        rom[327][52] = -8'd22;
        rom[327][53] = -8'd29;
        rom[327][54] = -8'd4;
        rom[327][55] = -8'd8;
        rom[327][56] = -8'd1;
        rom[327][57] = -8'd25;
        rom[327][58] = -8'd2;
        rom[327][59] = -8'd11;
        rom[327][60] = -8'd43;
        rom[327][61] = -8'd10;
        rom[327][62] = 8'd22;
        rom[327][63] = 8'd2;
        rom[328][0] = 8'd18;
        rom[328][1] = 8'd24;
        rom[328][2] = 8'd22;
        rom[328][3] = 8'd11;
        rom[328][4] = -8'd4;
        rom[328][5] = 8'd14;
        rom[328][6] = -8'd36;
        rom[328][7] = 8'd4;
        rom[328][8] = 8'd2;
        rom[328][9] = -8'd13;
        rom[328][10] = -8'd68;
        rom[328][11] = 8'd24;
        rom[328][12] = -8'd22;
        rom[328][13] = -8'd8;
        rom[328][14] = 8'd14;
        rom[328][15] = 8'd14;
        rom[328][16] = 8'd5;
        rom[328][17] = -8'd41;
        rom[328][18] = -8'd21;
        rom[328][19] = 8'd16;
        rom[328][20] = -8'd12;
        rom[328][21] = -8'd5;
        rom[328][22] = -8'd3;
        rom[328][23] = -8'd4;
        rom[328][24] = -8'd5;
        rom[328][25] = 8'd42;
        rom[328][26] = 8'd22;
        rom[328][27] = -8'd17;
        rom[328][28] = -8'd1;
        rom[328][29] = 8'd13;
        rom[328][30] = 8'd23;
        rom[328][31] = 8'd9;
        rom[328][32] = 8'd20;
        rom[328][33] = -8'd15;
        rom[328][34] = -8'd9;
        rom[328][35] = 8'd8;
        rom[328][36] = -8'd11;
        rom[328][37] = 8'd12;
        rom[328][38] = -8'd63;
        rom[328][39] = -8'd13;
        rom[328][40] = -8'd10;
        rom[328][41] = -8'd32;
        rom[328][42] = -8'd5;
        rom[328][43] = 8'd8;
        rom[328][44] = 8'd35;
        rom[328][45] = -8'd9;
        rom[328][46] = 8'd16;
        rom[328][47] = 8'd26;
        rom[328][48] = 8'd3;
        rom[328][49] = 8'd10;
        rom[328][50] = 8'd6;
        rom[328][51] = 8'd7;
        rom[328][52] = -8'd6;
        rom[328][53] = -8'd4;
        rom[328][54] = -8'd7;
        rom[328][55] = 8'd4;
        rom[328][56] = -8'd23;
        rom[328][57] = 8'd3;
        rom[328][58] = 8'd10;
        rom[328][59] = -8'd26;
        rom[328][60] = -8'd9;
        rom[328][61] = -8'd11;
        rom[328][62] = -8'd5;
        rom[328][63] = -8'd36;
        rom[329][0] = -8'd25;
        rom[329][1] = -8'd17;
        rom[329][2] = 8'd5;
        rom[329][3] = 8'd32;
        rom[329][4] = -8'd22;
        rom[329][5] = 8'd1;
        rom[329][6] = -8'd38;
        rom[329][7] = -8'd11;
        rom[329][8] = 8'd15;
        rom[329][9] = -8'd1;
        rom[329][10] = -8'd15;
        rom[329][11] = 8'd38;
        rom[329][12] = 8'd11;
        rom[329][13] = 8'd14;
        rom[329][14] = 8'd16;
        rom[329][15] = 8'd5;
        rom[329][16] = -8'd7;
        rom[329][17] = 8'd24;
        rom[329][18] = 8'd57;
        rom[329][19] = -8'd33;
        rom[329][20] = 8'd6;
        rom[329][21] = 8'd4;
        rom[329][22] = 8'd7;
        rom[329][23] = -8'd6;
        rom[329][24] = 8'd5;
        rom[329][25] = 8'd0;
        rom[329][26] = 8'd6;
        rom[329][27] = -8'd8;
        rom[329][28] = -8'd33;
        rom[329][29] = -8'd18;
        rom[329][30] = -8'd1;
        rom[329][31] = 8'd20;
        rom[329][32] = 8'd2;
        rom[329][33] = -8'd17;
        rom[329][34] = 8'd41;
        rom[329][35] = 8'd21;
        rom[329][36] = 8'd8;
        rom[329][37] = -8'd7;
        rom[329][38] = 8'd5;
        rom[329][39] = -8'd28;
        rom[329][40] = -8'd11;
        rom[329][41] = -8'd4;
        rom[329][42] = 8'd41;
        rom[329][43] = 8'd13;
        rom[329][44] = -8'd7;
        rom[329][45] = -8'd9;
        rom[329][46] = -8'd13;
        rom[329][47] = 8'd22;
        rom[329][48] = 8'd0;
        rom[329][49] = -8'd24;
        rom[329][50] = 8'd26;
        rom[329][51] = 8'd31;
        rom[329][52] = 8'd6;
        rom[329][53] = 8'd12;
        rom[329][54] = 8'd9;
        rom[329][55] = 8'd7;
        rom[329][56] = -8'd38;
        rom[329][57] = -8'd19;
        rom[329][58] = -8'd3;
        rom[329][59] = 8'd62;
        rom[329][60] = -8'd33;
        rom[329][61] = 8'd31;
        rom[329][62] = -8'd28;
        rom[329][63] = 8'd9;
        rom[330][0] = 8'd24;
        rom[330][1] = -8'd24;
        rom[330][2] = 8'd33;
        rom[330][3] = -8'd36;
        rom[330][4] = -8'd5;
        rom[330][5] = -8'd3;
        rom[330][6] = -8'd8;
        rom[330][7] = -8'd5;
        rom[330][8] = -8'd1;
        rom[330][9] = 8'd17;
        rom[330][10] = -8'd35;
        rom[330][11] = -8'd21;
        rom[330][12] = 8'd28;
        rom[330][13] = -8'd1;
        rom[330][14] = 8'd20;
        rom[330][15] = 8'd31;
        rom[330][16] = -8'd52;
        rom[330][17] = 8'd11;
        rom[330][18] = 8'd19;
        rom[330][19] = 8'd4;
        rom[330][20] = 8'd0;
        rom[330][21] = -8'd4;
        rom[330][22] = -8'd6;
        rom[330][23] = -8'd8;
        rom[330][24] = -8'd2;
        rom[330][25] = -8'd6;
        rom[330][26] = -8'd53;
        rom[330][27] = 8'd13;
        rom[330][28] = 8'd3;
        rom[330][29] = -8'd25;
        rom[330][30] = -8'd3;
        rom[330][31] = 8'd7;
        rom[330][32] = 8'd14;
        rom[330][33] = 8'd16;
        rom[330][34] = 8'd19;
        rom[330][35] = -8'd38;
        rom[330][36] = 8'd4;
        rom[330][37] = 8'd7;
        rom[330][38] = 8'd20;
        rom[330][39] = 8'd16;
        rom[330][40] = 8'd8;
        rom[330][41] = 8'd56;
        rom[330][42] = -8'd29;
        rom[330][43] = 8'd8;
        rom[330][44] = 8'd9;
        rom[330][45] = 8'd15;
        rom[330][46] = -8'd8;
        rom[330][47] = -8'd27;
        rom[330][48] = -8'd3;
        rom[330][49] = 8'd5;
        rom[330][50] = 8'd41;
        rom[330][51] = -8'd17;
        rom[330][52] = 8'd12;
        rom[330][53] = 8'd21;
        rom[330][54] = 8'd23;
        rom[330][55] = -8'd26;
        rom[330][56] = -8'd44;
        rom[330][57] = 8'd9;
        rom[330][58] = -8'd3;
        rom[330][59] = -8'd19;
        rom[330][60] = 8'd12;
        rom[330][61] = -8'd6;
        rom[330][62] = -8'd40;
        rom[330][63] = 8'd11;
        rom[331][0] = -8'd29;
        rom[331][1] = -8'd24;
        rom[331][2] = 8'd2;
        rom[331][3] = -8'd19;
        rom[331][4] = -8'd19;
        rom[331][5] = 8'd10;
        rom[331][6] = -8'd12;
        rom[331][7] = -8'd37;
        rom[331][8] = -8'd26;
        rom[331][9] = 8'd8;
        rom[331][10] = 8'd35;
        rom[331][11] = 8'd24;
        rom[331][12] = -8'd27;
        rom[331][13] = -8'd32;
        rom[331][14] = 8'd27;
        rom[331][15] = 8'd32;
        rom[331][16] = 8'd13;
        rom[331][17] = -8'd32;
        rom[331][18] = -8'd57;
        rom[331][19] = -8'd1;
        rom[331][20] = -8'd6;
        rom[331][21] = 8'd31;
        rom[331][22] = -8'd2;
        rom[331][23] = -8'd11;
        rom[331][24] = 8'd10;
        rom[331][25] = -8'd11;
        rom[331][26] = 8'd23;
        rom[331][27] = -8'd37;
        rom[331][28] = 8'd76;
        rom[331][29] = 8'd29;
        rom[331][30] = 8'd46;
        rom[331][31] = -8'd83;
        rom[331][32] = -8'd32;
        rom[331][33] = 8'd14;
        rom[331][34] = 8'd47;
        rom[331][35] = -8'd36;
        rom[331][36] = -8'd39;
        rom[331][37] = -8'd33;
        rom[331][38] = 8'd22;
        rom[331][39] = 8'd2;
        rom[331][40] = -8'd13;
        rom[331][41] = -8'd58;
        rom[331][42] = 8'd0;
        rom[331][43] = -8'd18;
        rom[331][44] = -8'd62;
        rom[331][45] = -8'd33;
        rom[331][46] = 8'd41;
        rom[331][47] = -8'd44;
        rom[331][48] = 8'd34;
        rom[331][49] = -8'd68;
        rom[331][50] = -8'd22;
        rom[331][51] = 8'd2;
        rom[331][52] = -8'd23;
        rom[331][53] = -8'd30;
        rom[331][54] = -8'd11;
        rom[331][55] = -8'd21;
        rom[331][56] = -8'd17;
        rom[331][57] = 8'd13;
        rom[331][58] = 8'd18;
        rom[331][59] = 8'd46;
        rom[331][60] = -8'd41;
        rom[331][61] = -8'd27;
        rom[331][62] = 8'd16;
        rom[331][63] = 8'd25;
        rom[332][0] = -8'd7;
        rom[332][1] = -8'd36;
        rom[332][2] = 8'd38;
        rom[332][3] = 8'd12;
        rom[332][4] = 8'd42;
        rom[332][5] = 8'd3;
        rom[332][6] = -8'd30;
        rom[332][7] = -8'd48;
        rom[332][8] = 8'd28;
        rom[332][9] = 8'd24;
        rom[332][10] = -8'd25;
        rom[332][11] = -8'd38;
        rom[332][12] = 8'd2;
        rom[332][13] = -8'd1;
        rom[332][14] = 8'd29;
        rom[332][15] = 8'd16;
        rom[332][16] = -8'd13;
        rom[332][17] = 8'd15;
        rom[332][18] = 8'd19;
        rom[332][19] = -8'd55;
        rom[332][20] = -8'd5;
        rom[332][21] = 8'd10;
        rom[332][22] = -8'd2;
        rom[332][23] = 8'd13;
        rom[332][24] = -8'd4;
        rom[332][25] = 8'd20;
        rom[332][26] = -8'd24;
        rom[332][27] = 8'd6;
        rom[332][28] = 8'd16;
        rom[332][29] = 8'd2;
        rom[332][30] = -8'd30;
        rom[332][31] = 8'd39;
        rom[332][32] = 8'd10;
        rom[332][33] = 8'd6;
        rom[332][34] = -8'd26;
        rom[332][35] = 8'd21;
        rom[332][36] = 8'd15;
        rom[332][37] = -8'd13;
        rom[332][38] = 8'd18;
        rom[332][39] = -8'd1;
        rom[332][40] = -8'd29;
        rom[332][41] = 8'd9;
        rom[332][42] = 8'd4;
        rom[332][43] = 8'd2;
        rom[332][44] = 8'd20;
        rom[332][45] = 8'd21;
        rom[332][46] = -8'd36;
        rom[332][47] = 8'd76;
        rom[332][48] = 8'd16;
        rom[332][49] = 8'd2;
        rom[332][50] = 8'd33;
        rom[332][51] = -8'd15;
        rom[332][52] = -8'd34;
        rom[332][53] = 8'd6;
        rom[332][54] = 8'd8;
        rom[332][55] = 8'd3;
        rom[332][56] = 8'd36;
        rom[332][57] = 8'd47;
        rom[332][58] = -8'd6;
        rom[332][59] = -8'd26;
        rom[332][60] = -8'd3;
        rom[332][61] = 8'd0;
        rom[332][62] = 8'd17;
        rom[332][63] = 8'd6;
        rom[333][0] = 8'd19;
        rom[333][1] = -8'd15;
        rom[333][2] = 8'd15;
        rom[333][3] = -8'd12;
        rom[333][4] = 8'd0;
        rom[333][5] = 8'd23;
        rom[333][6] = 8'd31;
        rom[333][7] = 8'd26;
        rom[333][8] = 8'd11;
        rom[333][9] = -8'd19;
        rom[333][10] = -8'd12;
        rom[333][11] = -8'd17;
        rom[333][12] = 8'd28;
        rom[333][13] = 8'd22;
        rom[333][14] = 8'd21;
        rom[333][15] = -8'd8;
        rom[333][16] = -8'd8;
        rom[333][17] = -8'd39;
        rom[333][18] = 8'd11;
        rom[333][19] = 8'd0;
        rom[333][20] = 8'd2;
        rom[333][21] = -8'd1;
        rom[333][22] = -8'd7;
        rom[333][23] = -8'd8;
        rom[333][24] = -8'd1;
        rom[333][25] = -8'd38;
        rom[333][26] = -8'd15;
        rom[333][27] = -8'd20;
        rom[333][28] = -8'd51;
        rom[333][29] = 8'd17;
        rom[333][30] = 8'd17;
        rom[333][31] = 8'd4;
        rom[333][32] = -8'd9;
        rom[333][33] = -8'd1;
        rom[333][34] = -8'd34;
        rom[333][35] = -8'd35;
        rom[333][36] = -8'd18;
        rom[333][37] = 8'd7;
        rom[333][38] = 8'd8;
        rom[333][39] = 8'd4;
        rom[333][40] = -8'd4;
        rom[333][41] = -8'd16;
        rom[333][42] = -8'd40;
        rom[333][43] = 8'd3;
        rom[333][44] = -8'd5;
        rom[333][45] = 8'd3;
        rom[333][46] = 8'd14;
        rom[333][47] = -8'd56;
        rom[333][48] = 8'd10;
        rom[333][49] = -8'd19;
        rom[333][50] = 8'd14;
        rom[333][51] = -8'd19;
        rom[333][52] = 8'd21;
        rom[333][53] = 8'd12;
        rom[333][54] = -8'd13;
        rom[333][55] = -8'd26;
        rom[333][56] = -8'd13;
        rom[333][57] = 8'd15;
        rom[333][58] = 8'd6;
        rom[333][59] = 8'd26;
        rom[333][60] = -8'd12;
        rom[333][61] = 8'd0;
        rom[333][62] = 8'd54;
        rom[333][63] = 8'd22;
        rom[334][0] = 8'd1;
        rom[334][1] = -8'd4;
        rom[334][2] = 8'd13;
        rom[334][3] = 8'd0;
        rom[334][4] = 8'd4;
        rom[334][5] = -8'd34;
        rom[334][6] = 8'd2;
        rom[334][7] = -8'd4;
        rom[334][8] = 8'd17;
        rom[334][9] = -8'd23;
        rom[334][10] = -8'd33;
        rom[334][11] = -8'd36;
        rom[334][12] = -8'd39;
        rom[334][13] = -8'd11;
        rom[334][14] = 8'd10;
        rom[334][15] = 8'd23;
        rom[334][16] = 8'd27;
        rom[334][17] = -8'd14;
        rom[334][18] = -8'd13;
        rom[334][19] = -8'd31;
        rom[334][20] = -8'd4;
        rom[334][21] = 8'd11;
        rom[334][22] = -8'd44;
        rom[334][23] = -8'd8;
        rom[334][24] = -8'd37;
        rom[334][25] = -8'd3;
        rom[334][26] = 8'd9;
        rom[334][27] = 8'd4;
        rom[334][28] = 8'd2;
        rom[334][29] = -8'd9;
        rom[334][30] = 8'd8;
        rom[334][31] = -8'd17;
        rom[334][32] = -8'd4;
        rom[334][33] = -8'd8;
        rom[334][34] = -8'd6;
        rom[334][35] = -8'd2;
        rom[334][36] = -8'd4;
        rom[334][37] = 8'd16;
        rom[334][38] = -8'd39;
        rom[334][39] = 8'd19;
        rom[334][40] = -8'd35;
        rom[334][41] = -8'd26;
        rom[334][42] = -8'd40;
        rom[334][43] = 8'd15;
        rom[334][44] = 8'd33;
        rom[334][45] = -8'd67;
        rom[334][46] = 8'd31;
        rom[334][47] = -8'd18;
        rom[334][48] = -8'd15;
        rom[334][49] = -8'd18;
        rom[334][50] = 8'd4;
        rom[334][51] = 8'd22;
        rom[334][52] = -8'd1;
        rom[334][53] = -8'd3;
        rom[334][54] = -8'd13;
        rom[334][55] = -8'd40;
        rom[334][56] = -8'd13;
        rom[334][57] = 8'd17;
        rom[334][58] = 8'd17;
        rom[334][59] = -8'd3;
        rom[334][60] = -8'd30;
        rom[334][61] = -8'd27;
        rom[334][62] = 8'd25;
        rom[334][63] = -8'd16;
        rom[335][0] = 8'd13;
        rom[335][1] = -8'd42;
        rom[335][2] = -8'd15;
        rom[335][3] = 8'd15;
        rom[335][4] = 8'd29;
        rom[335][5] = -8'd23;
        rom[335][6] = 8'd10;
        rom[335][7] = 8'd0;
        rom[335][8] = 8'd29;
        rom[335][9] = 8'd48;
        rom[335][10] = -8'd10;
        rom[335][11] = -8'd6;
        rom[335][12] = -8'd42;
        rom[335][13] = 8'd6;
        rom[335][14] = 8'd23;
        rom[335][15] = -8'd1;
        rom[335][16] = -8'd6;
        rom[335][17] = -8'd10;
        rom[335][18] = 8'd2;
        rom[335][19] = -8'd11;
        rom[335][20] = 8'd0;
        rom[335][21] = 8'd13;
        rom[335][22] = 8'd12;
        rom[335][23] = 8'd15;
        rom[335][24] = -8'd54;
        rom[335][25] = -8'd4;
        rom[335][26] = -8'd8;
        rom[335][27] = -8'd28;
        rom[335][28] = -8'd10;
        rom[335][29] = 8'd6;
        rom[335][30] = -8'd5;
        rom[335][31] = 8'd15;
        rom[335][32] = -8'd27;
        rom[335][33] = 8'd14;
        rom[335][34] = 8'd16;
        rom[335][35] = 8'd35;
        rom[335][36] = -8'd17;
        rom[335][37] = -8'd3;
        rom[335][38] = 8'd11;
        rom[335][39] = -8'd10;
        rom[335][40] = 8'd9;
        rom[335][41] = -8'd4;
        rom[335][42] = 8'd3;
        rom[335][43] = -8'd37;
        rom[335][44] = 8'd1;
        rom[335][45] = -8'd24;
        rom[335][46] = -8'd6;
        rom[335][47] = 8'd13;
        rom[335][48] = 8'd20;
        rom[335][49] = -8'd16;
        rom[335][50] = -8'd49;
        rom[335][51] = 8'd15;
        rom[335][52] = 8'd10;
        rom[335][53] = 8'd29;
        rom[335][54] = -8'd32;
        rom[335][55] = -8'd44;
        rom[335][56] = 8'd23;
        rom[335][57] = -8'd26;
        rom[335][58] = -8'd24;
        rom[335][59] = 8'd0;
        rom[335][60] = 8'd48;
        rom[335][61] = -8'd23;
        rom[335][62] = -8'd29;
        rom[335][63] = -8'd9;
        rom[336][0] = 8'd8;
        rom[336][1] = 8'd0;
        rom[336][2] = -8'd2;
        rom[336][3] = 8'd10;
        rom[336][4] = -8'd8;
        rom[336][5] = -8'd2;
        rom[336][6] = 8'd2;
        rom[336][7] = 8'd6;
        rom[336][8] = 8'd0;
        rom[336][9] = -8'd1;
        rom[336][10] = -8'd6;
        rom[336][11] = -8'd10;
        rom[336][12] = 8'd7;
        rom[336][13] = 8'd4;
        rom[336][14] = 8'd4;
        rom[336][15] = 8'd8;
        rom[336][16] = 8'd8;
        rom[336][17] = -8'd5;
        rom[336][18] = -8'd5;
        rom[336][19] = 8'd0;
        rom[336][20] = -8'd2;
        rom[336][21] = 8'd0;
        rom[336][22] = 8'd3;
        rom[336][23] = 8'd4;
        rom[336][24] = -8'd6;
        rom[336][25] = -8'd8;
        rom[336][26] = 8'd2;
        rom[336][27] = -8'd4;
        rom[336][28] = 8'd7;
        rom[336][29] = -8'd8;
        rom[336][30] = 8'd5;
        rom[336][31] = 8'd0;
        rom[336][32] = 8'd4;
        rom[336][33] = -8'd4;
        rom[336][34] = 8'd7;
        rom[336][35] = -8'd6;
        rom[336][36] = 8'd3;
        rom[336][37] = -8'd6;
        rom[336][38] = -8'd6;
        rom[336][39] = 8'd7;
        rom[336][40] = -8'd2;
        rom[336][41] = 8'd1;
        rom[336][42] = 8'd1;
        rom[336][43] = -8'd6;
        rom[336][44] = -8'd3;
        rom[336][45] = 8'd0;
        rom[336][46] = 8'd1;
        rom[336][47] = -8'd2;
        rom[336][48] = 8'd9;
        rom[336][49] = 8'd1;
        rom[336][50] = 8'd2;
        rom[336][51] = -8'd7;
        rom[336][52] = -8'd1;
        rom[336][53] = 8'd7;
        rom[336][54] = 8'd3;
        rom[336][55] = 8'd4;
        rom[336][56] = -8'd5;
        rom[336][57] = 8'd9;
        rom[336][58] = 8'd4;
        rom[336][59] = 8'd3;
        rom[336][60] = -8'd1;
        rom[336][61] = -8'd1;
        rom[336][62] = 8'd0;
        rom[336][63] = -8'd1;
        rom[337][0] = -8'd14;
        rom[337][1] = 8'd30;
        rom[337][2] = -8'd76;
        rom[337][3] = 8'd30;
        rom[337][4] = -8'd29;
        rom[337][5] = -8'd47;
        rom[337][6] = 8'd18;
        rom[337][7] = 8'd19;
        rom[337][8] = 8'd0;
        rom[337][9] = -8'd5;
        rom[337][10] = -8'd19;
        rom[337][11] = -8'd4;
        rom[337][12] = 8'd13;
        rom[337][13] = -8'd2;
        rom[337][14] = -8'd19;
        rom[337][15] = 8'd12;
        rom[337][16] = 8'd16;
        rom[337][17] = -8'd6;
        rom[337][18] = 8'd0;
        rom[337][19] = -8'd33;
        rom[337][20] = -8'd4;
        rom[337][21] = 8'd8;
        rom[337][22] = -8'd51;
        rom[337][23] = -8'd111;
        rom[337][24] = -8'd30;
        rom[337][25] = 8'd11;
        rom[337][26] = -8'd5;
        rom[337][27] = -8'd66;
        rom[337][28] = 8'd23;
        rom[337][29] = 8'd14;
        rom[337][30] = -8'd3;
        rom[337][31] = 8'd21;
        rom[337][32] = 8'd15;
        rom[337][33] = 8'd13;
        rom[337][34] = 8'd0;
        rom[337][35] = -8'd24;
        rom[337][36] = -8'd19;
        rom[337][37] = 8'd30;
        rom[337][38] = -8'd1;
        rom[337][39] = -8'd1;
        rom[337][40] = -8'd7;
        rom[337][41] = -8'd13;
        rom[337][42] = 8'd2;
        rom[337][43] = 8'd24;
        rom[337][44] = -8'd4;
        rom[337][45] = -8'd12;
        rom[337][46] = 8'd6;
        rom[337][47] = -8'd11;
        rom[337][48] = -8'd30;
        rom[337][49] = 8'd7;
        rom[337][50] = -8'd18;
        rom[337][51] = 8'd64;
        rom[337][52] = 8'd21;
        rom[337][53] = 8'd17;
        rom[337][54] = -8'd3;
        rom[337][55] = 8'd61;
        rom[337][56] = -8'd10;
        rom[337][57] = -8'd11;
        rom[337][58] = -8'd12;
        rom[337][59] = 8'd3;
        rom[337][60] = 8'd27;
        rom[337][61] = -8'd4;
        rom[337][62] = -8'd34;
        rom[337][63] = -8'd15;
        rom[338][0] = 8'd0;
        rom[338][1] = 8'd32;
        rom[338][2] = 8'd29;
        rom[338][3] = -8'd21;
        rom[338][4] = -8'd21;
        rom[338][5] = 8'd6;
        rom[338][6] = 8'd4;
        rom[338][7] = 8'd3;
        rom[338][8] = 8'd20;
        rom[338][9] = 8'd3;
        rom[338][10] = -8'd20;
        rom[338][11] = 8'd11;
        rom[338][12] = 8'd5;
        rom[338][13] = -8'd32;
        rom[338][14] = 8'd35;
        rom[338][15] = -8'd1;
        rom[338][16] = -8'd51;
        rom[338][17] = 8'd8;
        rom[338][18] = 8'd10;
        rom[338][19] = 8'd2;
        rom[338][20] = -8'd13;
        rom[338][21] = 8'd2;
        rom[338][22] = -8'd3;
        rom[338][23] = -8'd26;
        rom[338][24] = -8'd8;
        rom[338][25] = 8'd2;
        rom[338][26] = 8'd34;
        rom[338][27] = -8'd8;
        rom[338][28] = -8'd14;
        rom[338][29] = -8'd13;
        rom[338][30] = 8'd9;
        rom[338][31] = -8'd6;
        rom[338][32] = -8'd25;
        rom[338][33] = 8'd11;
        rom[338][34] = -8'd4;
        rom[338][35] = 8'd3;
        rom[338][36] = -8'd25;
        rom[338][37] = -8'd3;
        rom[338][38] = 8'd7;
        rom[338][39] = -8'd6;
        rom[338][40] = 8'd4;
        rom[338][41] = 8'd5;
        rom[338][42] = 8'd5;
        rom[338][43] = -8'd8;
        rom[338][44] = -8'd24;
        rom[338][45] = -8'd4;
        rom[338][46] = -8'd25;
        rom[338][47] = -8'd31;
        rom[338][48] = 8'd25;
        rom[338][49] = -8'd21;
        rom[338][50] = 8'd0;
        rom[338][51] = 8'd21;
        rom[338][52] = -8'd26;
        rom[338][53] = 8'd21;
        rom[338][54] = 8'd21;
        rom[338][55] = 8'd10;
        rom[338][56] = 8'd5;
        rom[338][57] = 8'd19;
        rom[338][58] = -8'd68;
        rom[338][59] = -8'd10;
        rom[338][60] = -8'd12;
        rom[338][61] = -8'd34;
        rom[338][62] = -8'd2;
        rom[338][63] = -8'd6;
        rom[339][0] = 8'd5;
        rom[339][1] = -8'd80;
        rom[339][2] = -8'd48;
        rom[339][3] = -8'd40;
        rom[339][4] = 8'd8;
        rom[339][5] = -8'd6;
        rom[339][6] = -8'd56;
        rom[339][7] = -8'd20;
        rom[339][8] = -8'd56;
        rom[339][9] = 8'd2;
        rom[339][10] = -8'd72;
        rom[339][11] = -8'd25;
        rom[339][12] = 8'd15;
        rom[339][13] = 8'd21;
        rom[339][14] = 8'd33;
        rom[339][15] = -8'd8;
        rom[339][16] = 8'd7;
        rom[339][17] = -8'd31;
        rom[339][18] = -8'd16;
        rom[339][19] = -8'd12;
        rom[339][20] = -8'd4;
        rom[339][21] = -8'd6;
        rom[339][22] = -8'd29;
        rom[339][23] = -8'd12;
        rom[339][24] = 8'd1;
        rom[339][25] = 8'd8;
        rom[339][26] = 8'd15;
        rom[339][27] = -8'd1;
        rom[339][28] = 8'd14;
        rom[339][29] = -8'd30;
        rom[339][30] = -8'd29;
        rom[339][31] = 8'd12;
        rom[339][32] = -8'd17;
        rom[339][33] = 8'd26;
        rom[339][34] = 8'd23;
        rom[339][35] = -8'd4;
        rom[339][36] = 8'd1;
        rom[339][37] = 8'd5;
        rom[339][38] = 8'd21;
        rom[339][39] = -8'd25;
        rom[339][40] = -8'd9;
        rom[339][41] = 8'd19;
        rom[339][42] = -8'd18;
        rom[339][43] = -8'd67;
        rom[339][44] = -8'd9;
        rom[339][45] = 8'd4;
        rom[339][46] = 8'd22;
        rom[339][47] = 8'd25;
        rom[339][48] = 8'd23;
        rom[339][49] = 8'd11;
        rom[339][50] = 8'd12;
        rom[339][51] = 8'd31;
        rom[339][52] = 8'd21;
        rom[339][53] = -8'd3;
        rom[339][54] = -8'd51;
        rom[339][55] = -8'd17;
        rom[339][56] = -8'd11;
        rom[339][57] = 8'd15;
        rom[339][58] = 8'd3;
        rom[339][59] = -8'd9;
        rom[339][60] = -8'd2;
        rom[339][61] = -8'd17;
        rom[339][62] = -8'd2;
        rom[339][63] = -8'd12;
        rom[340][0] = 8'd9;
        rom[340][1] = 8'd28;
        rom[340][2] = -8'd22;
        rom[340][3] = 8'd3;
        rom[340][4] = -8'd18;
        rom[340][5] = -8'd5;
        rom[340][6] = 8'd30;
        rom[340][7] = -8'd29;
        rom[340][8] = 8'd9;
        rom[340][9] = 8'd3;
        rom[340][10] = -8'd19;
        rom[340][11] = -8'd6;
        rom[340][12] = -8'd19;
        rom[340][13] = -8'd65;
        rom[340][14] = -8'd52;
        rom[340][15] = -8'd36;
        rom[340][16] = 8'd19;
        rom[340][17] = 8'd16;
        rom[340][18] = -8'd12;
        rom[340][19] = -8'd12;
        rom[340][20] = 8'd0;
        rom[340][21] = -8'd23;
        rom[340][22] = 8'd1;
        rom[340][23] = 8'd8;
        rom[340][24] = -8'd12;
        rom[340][25] = -8'd33;
        rom[340][26] = -8'd7;
        rom[340][27] = -8'd25;
        rom[340][28] = -8'd31;
        rom[340][29] = -8'd4;
        rom[340][30] = -8'd40;
        rom[340][31] = -8'd3;
        rom[340][32] = -8'd47;
        rom[340][33] = -8'd7;
        rom[340][34] = -8'd7;
        rom[340][35] = -8'd1;
        rom[340][36] = -8'd9;
        rom[340][37] = 8'd10;
        rom[340][38] = 8'd31;
        rom[340][39] = -8'd22;
        rom[340][40] = 8'd9;
        rom[340][41] = 8'd24;
        rom[340][42] = 8'd27;
        rom[340][43] = -8'd32;
        rom[340][44] = -8'd16;
        rom[340][45] = 8'd7;
        rom[340][46] = -8'd9;
        rom[340][47] = 8'd60;
        rom[340][48] = -8'd13;
        rom[340][49] = 8'd14;
        rom[340][50] = -8'd20;
        rom[340][51] = 8'd9;
        rom[340][52] = -8'd41;
        rom[340][53] = -8'd2;
        rom[340][54] = 8'd3;
        rom[340][55] = 8'd18;
        rom[340][56] = -8'd38;
        rom[340][57] = -8'd9;
        rom[340][58] = 8'd36;
        rom[340][59] = -8'd2;
        rom[340][60] = -8'd1;
        rom[340][61] = -8'd51;
        rom[340][62] = -8'd24;
        rom[340][63] = 8'd5;
        rom[341][0] = -8'd3;
        rom[341][1] = 8'd5;
        rom[341][2] = 8'd4;
        rom[341][3] = 8'd1;
        rom[341][4] = 8'd1;
        rom[341][5] = -8'd6;
        rom[341][6] = -8'd9;
        rom[341][7] = 8'd0;
        rom[341][8] = 8'd11;
        rom[341][9] = -8'd3;
        rom[341][10] = -8'd4;
        rom[341][11] = -8'd8;
        rom[341][12] = -8'd1;
        rom[341][13] = 8'd9;
        rom[341][14] = -8'd1;
        rom[341][15] = 8'd2;
        rom[341][16] = -8'd3;
        rom[341][17] = 8'd6;
        rom[341][18] = -8'd4;
        rom[341][19] = -8'd4;
        rom[341][20] = 8'd4;
        rom[341][21] = 8'd4;
        rom[341][22] = -8'd1;
        rom[341][23] = -8'd4;
        rom[341][24] = -8'd2;
        rom[341][25] = -8'd7;
        rom[341][26] = -8'd3;
        rom[341][27] = 8'd7;
        rom[341][28] = -8'd6;
        rom[341][29] = -8'd2;
        rom[341][30] = 8'd8;
        rom[341][31] = 8'd2;
        rom[341][32] = 8'd1;
        rom[341][33] = -8'd5;
        rom[341][34] = 8'd0;
        rom[341][35] = -8'd10;
        rom[341][36] = -8'd6;
        rom[341][37] = -8'd4;
        rom[341][38] = 8'd3;
        rom[341][39] = 8'd5;
        rom[341][40] = 8'd7;
        rom[341][41] = 8'd8;
        rom[341][42] = 8'd7;
        rom[341][43] = -8'd3;
        rom[341][44] = 8'd4;
        rom[341][45] = 8'd9;
        rom[341][46] = -8'd1;
        rom[341][47] = -8'd4;
        rom[341][48] = 8'd0;
        rom[341][49] = -8'd8;
        rom[341][50] = 8'd5;
        rom[341][51] = 8'd3;
        rom[341][52] = 8'd0;
        rom[341][53] = -8'd11;
        rom[341][54] = -8'd5;
        rom[341][55] = -8'd9;
        rom[341][56] = -8'd1;
        rom[341][57] = -8'd1;
        rom[341][58] = -8'd6;
        rom[341][59] = -8'd2;
        rom[341][60] = -8'd5;
        rom[341][61] = -8'd8;
        rom[341][62] = 8'd5;
        rom[341][63] = 8'd2;
        rom[342][0] = -8'd29;
        rom[342][1] = 8'd26;
        rom[342][2] = -8'd23;
        rom[342][3] = -8'd10;
        rom[342][4] = -8'd62;
        rom[342][5] = -8'd102;
        rom[342][6] = -8'd8;
        rom[342][7] = -8'd5;
        rom[342][8] = -8'd22;
        rom[342][9] = 8'd7;
        rom[342][10] = -8'd31;
        rom[342][11] = 8'd13;
        rom[342][12] = -8'd39;
        rom[342][13] = -8'd24;
        rom[342][14] = -8'd10;
        rom[342][15] = 8'd10;
        rom[342][16] = 8'd48;
        rom[342][17] = 8'd20;
        rom[342][18] = -8'd41;
        rom[342][19] = 8'd13;
        rom[342][20] = -8'd4;
        rom[342][21] = 8'd12;
        rom[342][22] = -8'd15;
        rom[342][23] = -8'd51;
        rom[342][24] = 8'd4;
        rom[342][25] = 8'd36;
        rom[342][26] = -8'd34;
        rom[342][27] = -8'd29;
        rom[342][28] = 8'd6;
        rom[342][29] = -8'd22;
        rom[342][30] = -8'd11;
        rom[342][31] = -8'd12;
        rom[342][32] = -8'd60;
        rom[342][33] = 8'd38;
        rom[342][34] = 8'd9;
        rom[342][35] = -8'd74;
        rom[342][36] = 8'd32;
        rom[342][37] = 8'd49;
        rom[342][38] = 8'd33;
        rom[342][39] = -8'd2;
        rom[342][40] = -8'd68;
        rom[342][41] = 8'd0;
        rom[342][42] = 8'd10;
        rom[342][43] = -8'd9;
        rom[342][44] = -8'd5;
        rom[342][45] = -8'd7;
        rom[342][46] = 8'd22;
        rom[342][47] = -8'd101;
        rom[342][48] = 8'd17;
        rom[342][49] = -8'd36;
        rom[342][50] = -8'd24;
        rom[342][51] = -8'd19;
        rom[342][52] = 8'd27;
        rom[342][53] = 8'd10;
        rom[342][54] = 8'd19;
        rom[342][55] = -8'd38;
        rom[342][56] = -8'd3;
        rom[342][57] = -8'd29;
        rom[342][58] = -8'd64;
        rom[342][59] = 8'd27;
        rom[342][60] = -8'd37;
        rom[342][61] = -8'd17;
        rom[342][62] = 8'd10;
        rom[342][63] = 8'd9;
        rom[343][0] = 8'd2;
        rom[343][1] = 8'd5;
        rom[343][2] = -8'd17;
        rom[343][3] = -8'd5;
        rom[343][4] = 8'd5;
        rom[343][5] = 8'd35;
        rom[343][6] = -8'd9;
        rom[343][7] = -8'd23;
        rom[343][8] = -8'd40;
        rom[343][9] = -8'd3;
        rom[343][10] = -8'd15;
        rom[343][11] = 8'd8;
        rom[343][12] = 8'd14;
        rom[343][13] = 8'd48;
        rom[343][14] = -8'd6;
        rom[343][15] = -8'd42;
        rom[343][16] = -8'd23;
        rom[343][17] = -8'd13;
        rom[343][18] = -8'd6;
        rom[343][19] = 8'd15;
        rom[343][20] = 8'd1;
        rom[343][21] = -8'd7;
        rom[343][22] = -8'd12;
        rom[343][23] = -8'd11;
        rom[343][24] = 8'd19;
        rom[343][25] = -8'd13;
        rom[343][26] = -8'd42;
        rom[343][27] = 8'd6;
        rom[343][28] = -8'd19;
        rom[343][29] = 8'd15;
        rom[343][30] = 8'd17;
        rom[343][31] = 8'd26;
        rom[343][32] = -8'd4;
        rom[343][33] = -8'd19;
        rom[343][34] = 8'd3;
        rom[343][35] = -8'd5;
        rom[343][36] = -8'd9;
        rom[343][37] = -8'd1;
        rom[343][38] = 8'd26;
        rom[343][39] = 8'd9;
        rom[343][40] = 8'd27;
        rom[343][41] = -8'd1;
        rom[343][42] = -8'd7;
        rom[343][43] = 8'd11;
        rom[343][44] = -8'd4;
        rom[343][45] = -8'd10;
        rom[343][46] = -8'd18;
        rom[343][47] = 8'd50;
        rom[343][48] = -8'd28;
        rom[343][49] = 8'd21;
        rom[343][50] = 8'd7;
        rom[343][51] = 8'd0;
        rom[343][52] = -8'd2;
        rom[343][53] = -8'd28;
        rom[343][54] = -8'd4;
        rom[343][55] = -8'd17;
        rom[343][56] = -8'd14;
        rom[343][57] = -8'd28;
        rom[343][58] = -8'd6;
        rom[343][59] = -8'd31;
        rom[343][60] = 8'd4;
        rom[343][61] = -8'd11;
        rom[343][62] = 8'd21;
        rom[343][63] = 8'd25;
        rom[344][0] = -8'd13;
        rom[344][1] = 8'd4;
        rom[344][2] = -8'd12;
        rom[344][3] = 8'd11;
        rom[344][4] = -8'd22;
        rom[344][5] = -8'd1;
        rom[344][6] = -8'd35;
        rom[344][7] = 8'd27;
        rom[344][8] = -8'd10;
        rom[344][9] = -8'd30;
        rom[344][10] = -8'd11;
        rom[344][11] = 8'd4;
        rom[344][12] = 8'd20;
        rom[344][13] = 8'd26;
        rom[344][14] = -8'd4;
        rom[344][15] = 8'd27;
        rom[344][16] = 8'd12;
        rom[344][17] = -8'd2;
        rom[344][18] = -8'd16;
        rom[344][19] = 8'd23;
        rom[344][20] = -8'd12;
        rom[344][21] = -8'd17;
        rom[344][22] = 8'd10;
        rom[344][23] = 8'd0;
        rom[344][24] = 8'd7;
        rom[344][25] = 8'd2;
        rom[344][26] = 8'd4;
        rom[344][27] = 8'd67;
        rom[344][28] = -8'd16;
        rom[344][29] = 8'd29;
        rom[344][30] = -8'd5;
        rom[344][31] = -8'd17;
        rom[344][32] = 8'd35;
        rom[344][33] = 8'd32;
        rom[344][34] = 8'd15;
        rom[344][35] = 8'd8;
        rom[344][36] = 8'd2;
        rom[344][37] = 8'd44;
        rom[344][38] = 8'd19;
        rom[344][39] = -8'd2;
        rom[344][40] = 8'd27;
        rom[344][41] = -8'd1;
        rom[344][42] = 8'd20;
        rom[344][43] = 8'd7;
        rom[344][44] = -8'd62;
        rom[344][45] = 8'd33;
        rom[344][46] = 8'd0;
        rom[344][47] = -8'd46;
        rom[344][48] = -8'd53;
        rom[344][49] = 8'd6;
        rom[344][50] = 8'd4;
        rom[344][51] = 8'd17;
        rom[344][52] = 8'd12;
        rom[344][53] = -8'd13;
        rom[344][54] = 8'd17;
        rom[344][55] = 8'd41;
        rom[344][56] = 8'd7;
        rom[344][57] = -8'd15;
        rom[344][58] = 8'd33;
        rom[344][59] = 8'd7;
        rom[344][60] = 8'd6;
        rom[344][61] = 8'd31;
        rom[344][62] = 8'd2;
        rom[344][63] = 8'd24;
        rom[345][0] = 8'd8;
        rom[345][1] = 8'd17;
        rom[345][2] = -8'd10;
        rom[345][3] = -8'd16;
        rom[345][4] = -8'd31;
        rom[345][5] = -8'd20;
        rom[345][6] = 8'd6;
        rom[345][7] = 8'd13;
        rom[345][8] = -8'd11;
        rom[345][9] = -8'd4;
        rom[345][10] = 8'd13;
        rom[345][11] = -8'd33;
        rom[345][12] = 8'd56;
        rom[345][13] = -8'd43;
        rom[345][14] = 8'd14;
        rom[345][15] = 8'd31;
        rom[345][16] = -8'd7;
        rom[345][17] = 8'd49;
        rom[345][18] = 8'd33;
        rom[345][19] = 8'd33;
        rom[345][20] = -8'd16;
        rom[345][21] = -8'd27;
        rom[345][22] = -8'd32;
        rom[345][23] = 8'd26;
        rom[345][24] = -8'd31;
        rom[345][25] = 8'd24;
        rom[345][26] = 8'd0;
        rom[345][27] = -8'd6;
        rom[345][28] = 8'd8;
        rom[345][29] = 8'd23;
        rom[345][30] = -8'd7;
        rom[345][31] = 8'd6;
        rom[345][32] = -8'd6;
        rom[345][33] = 8'd19;
        rom[345][34] = -8'd10;
        rom[345][35] = -8'd16;
        rom[345][36] = 8'd8;
        rom[345][37] = -8'd21;
        rom[345][38] = 8'd3;
        rom[345][39] = -8'd9;
        rom[345][40] = -8'd57;
        rom[345][41] = 8'd32;
        rom[345][42] = -8'd45;
        rom[345][43] = -8'd14;
        rom[345][44] = 8'd10;
        rom[345][45] = 8'd7;
        rom[345][46] = -8'd5;
        rom[345][47] = -8'd68;
        rom[345][48] = 8'd24;
        rom[345][49] = 8'd11;
        rom[345][50] = -8'd24;
        rom[345][51] = -8'd51;
        rom[345][52] = -8'd21;
        rom[345][53] = -8'd2;
        rom[345][54] = 8'd8;
        rom[345][55] = -8'd23;
        rom[345][56] = 8'd0;
        rom[345][57] = 8'd7;
        rom[345][58] = 8'd32;
        rom[345][59] = 8'd13;
        rom[345][60] = -8'd2;
        rom[345][61] = 8'd16;
        rom[345][62] = -8'd6;
        rom[345][63] = 8'd30;
        rom[346][0] = -8'd26;
        rom[346][1] = 8'd35;
        rom[346][2] = 8'd1;
        rom[346][3] = -8'd46;
        rom[346][4] = 8'd5;
        rom[346][5] = 8'd20;
        rom[346][6] = 8'd19;
        rom[346][7] = -8'd35;
        rom[346][8] = -8'd22;
        rom[346][9] = 8'd10;
        rom[346][10] = 8'd14;
        rom[346][11] = -8'd25;
        rom[346][12] = 8'd5;
        rom[346][13] = -8'd8;
        rom[346][14] = -8'd30;
        rom[346][15] = -8'd37;
        rom[346][16] = 8'd14;
        rom[346][17] = 8'd15;
        rom[346][18] = -8'd35;
        rom[346][19] = 8'd7;
        rom[346][20] = -8'd1;
        rom[346][21] = 8'd3;
        rom[346][22] = 8'd22;
        rom[346][23] = -8'd39;
        rom[346][24] = -8'd8;
        rom[346][25] = -8'd4;
        rom[346][26] = -8'd53;
        rom[346][27] = 8'd1;
        rom[346][28] = 8'd5;
        rom[346][29] = 8'd30;
        rom[346][30] = 8'd7;
        rom[346][31] = -8'd4;
        rom[346][32] = -8'd21;
        rom[346][33] = -8'd15;
        rom[346][34] = 8'd3;
        rom[346][35] = 8'd0;
        rom[346][36] = -8'd20;
        rom[346][37] = 8'd19;
        rom[346][38] = -8'd38;
        rom[346][39] = 8'd20;
        rom[346][40] = 8'd23;
        rom[346][41] = 8'd7;
        rom[346][42] = 8'd19;
        rom[346][43] = 8'd28;
        rom[346][44] = 8'd16;
        rom[346][45] = -8'd27;
        rom[346][46] = 8'd3;
        rom[346][47] = -8'd13;
        rom[346][48] = -8'd7;
        rom[346][49] = 8'd5;
        rom[346][50] = -8'd19;
        rom[346][51] = -8'd6;
        rom[346][52] = 8'd6;
        rom[346][53] = -8'd14;
        rom[346][54] = -8'd9;
        rom[346][55] = -8'd35;
        rom[346][56] = -8'd1;
        rom[346][57] = -8'd2;
        rom[346][58] = -8'd8;
        rom[346][59] = -8'd20;
        rom[346][60] = -8'd13;
        rom[346][61] = -8'd47;
        rom[346][62] = -8'd11;
        rom[346][63] = 8'd43;
        rom[347][0] = -8'd13;
        rom[347][1] = -8'd11;
        rom[347][2] = 8'd6;
        rom[347][3] = -8'd1;
        rom[347][4] = -8'd17;
        rom[347][5] = 8'd2;
        rom[347][6] = -8'd17;
        rom[347][7] = -8'd22;
        rom[347][8] = 8'd16;
        rom[347][9] = 8'd15;
        rom[347][10] = 8'd23;
        rom[347][11] = 8'd12;
        rom[347][12] = -8'd21;
        rom[347][13] = 8'd17;
        rom[347][14] = -8'd19;
        rom[347][15] = -8'd9;
        rom[347][16] = 8'd30;
        rom[347][17] = 8'd3;
        rom[347][18] = 8'd23;
        rom[347][19] = -8'd9;
        rom[347][20] = -8'd4;
        rom[347][21] = 8'd20;
        rom[347][22] = -8'd16;
        rom[347][23] = 8'd44;
        rom[347][24] = -8'd40;
        rom[347][25] = 8'd10;
        rom[347][26] = -8'd4;
        rom[347][27] = -8'd1;
        rom[347][28] = -8'd12;
        rom[347][29] = 8'd5;
        rom[347][30] = -8'd3;
        rom[347][31] = -8'd10;
        rom[347][32] = -8'd5;
        rom[347][33] = 8'd34;
        rom[347][34] = -8'd1;
        rom[347][35] = 8'd13;
        rom[347][36] = 8'd4;
        rom[347][37] = 8'd33;
        rom[347][38] = 8'd0;
        rom[347][39] = -8'd3;
        rom[347][40] = 8'd20;
        rom[347][41] = 8'd1;
        rom[347][42] = 8'd9;
        rom[347][43] = -8'd31;
        rom[347][44] = -8'd16;
        rom[347][45] = 8'd44;
        rom[347][46] = 8'd42;
        rom[347][47] = 8'd37;
        rom[347][48] = 8'd19;
        rom[347][49] = -8'd17;
        rom[347][50] = 8'd12;
        rom[347][51] = -8'd7;
        rom[347][52] = 8'd6;
        rom[347][53] = -8'd15;
        rom[347][54] = 8'd29;
        rom[347][55] = 8'd7;
        rom[347][56] = 8'd17;
        rom[347][57] = -8'd58;
        rom[347][58] = 8'd19;
        rom[347][59] = 8'd41;
        rom[347][60] = 8'd4;
        rom[347][61] = 8'd12;
        rom[347][62] = 8'd3;
        rom[347][63] = -8'd40;
        rom[348][0] = -8'd49;
        rom[348][1] = -8'd25;
        rom[348][2] = 8'd0;
        rom[348][3] = -8'd7;
        rom[348][4] = 8'd15;
        rom[348][5] = 8'd22;
        rom[348][6] = 8'd18;
        rom[348][7] = 8'd45;
        rom[348][8] = -8'd10;
        rom[348][9] = 8'd11;
        rom[348][10] = -8'd16;
        rom[348][11] = 8'd4;
        rom[348][12] = -8'd11;
        rom[348][13] = 8'd18;
        rom[348][14] = 8'd3;
        rom[348][15] = 8'd21;
        rom[348][16] = -8'd36;
        rom[348][17] = -8'd15;
        rom[348][18] = -8'd68;
        rom[348][19] = 8'd6;
        rom[348][20] = -8'd12;
        rom[348][21] = -8'd18;
        rom[348][22] = -8'd7;
        rom[348][23] = -8'd31;
        rom[348][24] = -8'd4;
        rom[348][25] = 8'd1;
        rom[348][26] = -8'd34;
        rom[348][27] = -8'd6;
        rom[348][28] = -8'd1;
        rom[348][29] = 8'd19;
        rom[348][30] = 8'd22;
        rom[348][31] = 8'd9;
        rom[348][32] = -8'd20;
        rom[348][33] = -8'd29;
        rom[348][34] = 8'd2;
        rom[348][35] = 8'd9;
        rom[348][36] = 8'd33;
        rom[348][37] = -8'd13;
        rom[348][38] = 8'd28;
        rom[348][39] = 8'd9;
        rom[348][40] = -8'd50;
        rom[348][41] = 8'd23;
        rom[348][42] = -8'd9;
        rom[348][43] = 8'd22;
        rom[348][44] = 8'd13;
        rom[348][45] = 8'd8;
        rom[348][46] = 8'd12;
        rom[348][47] = 8'd8;
        rom[348][48] = -8'd19;
        rom[348][49] = 8'd2;
        rom[348][50] = 8'd0;
        rom[348][51] = 8'd15;
        rom[348][52] = 8'd11;
        rom[348][53] = 8'd4;
        rom[348][54] = 8'd9;
        rom[348][55] = -8'd8;
        rom[348][56] = 8'd5;
        rom[348][57] = 8'd12;
        rom[348][58] = -8'd8;
        rom[348][59] = 8'd36;
        rom[348][60] = 8'd23;
        rom[348][61] = 8'd23;
        rom[348][62] = 8'd14;
        rom[348][63] = 8'd6;
        rom[349][0] = -8'd13;
        rom[349][1] = -8'd20;
        rom[349][2] = -8'd13;
        rom[349][3] = -8'd27;
        rom[349][4] = 8'd21;
        rom[349][5] = 8'd2;
        rom[349][6] = -8'd7;
        rom[349][7] = -8'd28;
        rom[349][8] = -8'd8;
        rom[349][9] = 8'd12;
        rom[349][10] = -8'd14;
        rom[349][11] = 8'd0;
        rom[349][12] = -8'd19;
        rom[349][13] = 8'd37;
        rom[349][14] = 8'd24;
        rom[349][15] = -8'd11;
        rom[349][16] = 8'd10;
        rom[349][17] = -8'd4;
        rom[349][18] = -8'd13;
        rom[349][19] = -8'd28;
        rom[349][20] = 8'd1;
        rom[349][21] = 8'd26;
        rom[349][22] = -8'd11;
        rom[349][23] = -8'd26;
        rom[349][24] = -8'd5;
        rom[349][25] = -8'd12;
        rom[349][26] = -8'd3;
        rom[349][27] = 8'd18;
        rom[349][28] = -8'd5;
        rom[349][29] = -8'd27;
        rom[349][30] = -8'd51;
        rom[349][31] = 8'd6;
        rom[349][32] = -8'd6;
        rom[349][33] = 8'd32;
        rom[349][34] = 8'd12;
        rom[349][35] = 8'd5;
        rom[349][36] = 8'd6;
        rom[349][37] = 8'd4;
        rom[349][38] = -8'd6;
        rom[349][39] = -8'd61;
        rom[349][40] = -8'd2;
        rom[349][41] = 8'd8;
        rom[349][42] = -8'd38;
        rom[349][43] = -8'd9;
        rom[349][44] = 8'd5;
        rom[349][45] = 8'd34;
        rom[349][46] = 8'd7;
        rom[349][47] = 8'd32;
        rom[349][48] = -8'd17;
        rom[349][49] = -8'd30;
        rom[349][50] = -8'd23;
        rom[349][51] = -8'd9;
        rom[349][52] = 8'd0;
        rom[349][53] = -8'd2;
        rom[349][54] = -8'd39;
        rom[349][55] = 8'd18;
        rom[349][56] = -8'd35;
        rom[349][57] = 8'd8;
        rom[349][58] = 8'd8;
        rom[349][59] = -8'd51;
        rom[349][60] = -8'd61;
        rom[349][61] = 8'd21;
        rom[349][62] = -8'd12;
        rom[349][63] = -8'd33;
        rom[350][0] = 8'd19;
        rom[350][1] = -8'd37;
        rom[350][2] = 8'd31;
        rom[350][3] = 8'd0;
        rom[350][4] = -8'd57;
        rom[350][5] = 8'd3;
        rom[350][6] = 8'd7;
        rom[350][7] = 8'd9;
        rom[350][8] = 8'd9;
        rom[350][9] = -8'd20;
        rom[350][10] = -8'd3;
        rom[350][11] = 8'd27;
        rom[350][12] = -8'd26;
        rom[350][13] = -8'd1;
        rom[350][14] = 8'd19;
        rom[350][15] = -8'd1;
        rom[350][16] = -8'd7;
        rom[350][17] = 8'd3;
        rom[350][18] = 8'd7;
        rom[350][19] = -8'd7;
        rom[350][20] = 8'd0;
        rom[350][21] = -8'd15;
        rom[350][22] = -8'd38;
        rom[350][23] = 8'd5;
        rom[350][24] = 8'd4;
        rom[350][25] = 8'd1;
        rom[350][26] = -8'd2;
        rom[350][27] = -8'd17;
        rom[350][28] = 8'd2;
        rom[350][29] = -8'd42;
        rom[350][30] = -8'd25;
        rom[350][31] = -8'd6;
        rom[350][32] = 8'd9;
        rom[350][33] = -8'd57;
        rom[350][34] = -8'd44;
        rom[350][35] = 8'd13;
        rom[350][36] = 8'd1;
        rom[350][37] = -8'd5;
        rom[350][38] = -8'd17;
        rom[350][39] = 8'd30;
        rom[350][40] = 8'd4;
        rom[350][41] = -8'd24;
        rom[350][42] = -8'd3;
        rom[350][43] = -8'd21;
        rom[350][44] = -8'd17;
        rom[350][45] = 8'd13;
        rom[350][46] = 8'd18;
        rom[350][47] = 8'd4;
        rom[350][48] = 8'd40;
        rom[350][49] = -8'd55;
        rom[350][50] = -8'd32;
        rom[350][51] = 8'd7;
        rom[350][52] = 8'd5;
        rom[350][53] = -8'd1;
        rom[350][54] = -8'd22;
        rom[350][55] = 8'd12;
        rom[350][56] = -8'd17;
        rom[350][57] = -8'd25;
        rom[350][58] = -8'd16;
        rom[350][59] = 8'd12;
        rom[350][60] = -8'd12;
        rom[350][61] = 8'd36;
        rom[350][62] = 8'd59;
        rom[350][63] = 8'd18;
        rom[351][0] = -8'd2;
        rom[351][1] = -8'd34;
        rom[351][2] = 8'd3;
        rom[351][3] = -8'd5;
        rom[351][4] = -8'd16;
        rom[351][5] = -8'd70;
        rom[351][6] = 8'd4;
        rom[351][7] = -8'd5;
        rom[351][8] = -8'd28;
        rom[351][9] = -8'd40;
        rom[351][10] = -8'd12;
        rom[351][11] = -8'd8;
        rom[351][12] = 8'd9;
        rom[351][13] = -8'd17;
        rom[351][14] = 8'd24;
        rom[351][15] = 8'd35;
        rom[351][16] = -8'd8;
        rom[351][17] = 8'd10;
        rom[351][18] = -8'd42;
        rom[351][19] = 8'd10;
        rom[351][20] = -8'd9;
        rom[351][21] = -8'd4;
        rom[351][22] = 8'd3;
        rom[351][23] = -8'd33;
        rom[351][24] = -8'd1;
        rom[351][25] = -8'd21;
        rom[351][26] = -8'd7;
        rom[351][27] = -8'd26;
        rom[351][28] = -8'd18;
        rom[351][29] = -8'd5;
        rom[351][30] = 8'd25;
        rom[351][31] = -8'd28;
        rom[351][32] = 8'd10;
        rom[351][33] = 8'd15;
        rom[351][34] = 8'd13;
        rom[351][35] = -8'd7;
        rom[351][36] = 8'd6;
        rom[351][37] = 8'd32;
        rom[351][38] = 8'd3;
        rom[351][39] = 8'd22;
        rom[351][40] = -8'd30;
        rom[351][41] = -8'd5;
        rom[351][42] = -8'd16;
        rom[351][43] = 8'd11;
        rom[351][44] = -8'd22;
        rom[351][45] = -8'd78;
        rom[351][46] = -8'd35;
        rom[351][47] = -8'd14;
        rom[351][48] = -8'd65;
        rom[351][49] = -8'd2;
        rom[351][50] = 8'd15;
        rom[351][51] = -8'd1;
        rom[351][52] = -8'd35;
        rom[351][53] = 8'd42;
        rom[351][54] = -8'd62;
        rom[351][55] = 8'd17;
        rom[351][56] = -8'd70;
        rom[351][57] = -8'd13;
        rom[351][58] = -8'd16;
        rom[351][59] = -8'd4;
        rom[351][60] = 8'd24;
        rom[351][61] = 8'd30;
        rom[351][62] = -8'd29;
        rom[351][63] = -8'd12;
        rom[352][0] = 8'd21;
        rom[352][1] = -8'd1;
        rom[352][2] = 8'd33;
        rom[352][3] = 8'd15;
        rom[352][4] = -8'd1;
        rom[352][5] = 8'd22;
        rom[352][6] = 8'd22;
        rom[352][7] = 8'd33;
        rom[352][8] = 8'd9;
        rom[352][9] = 8'd2;
        rom[352][10] = -8'd47;
        rom[352][11] = 8'd7;
        rom[352][12] = -8'd44;
        rom[352][13] = -8'd38;
        rom[352][14] = 8'd6;
        rom[352][15] = -8'd33;
        rom[352][16] = -8'd41;
        rom[352][17] = 8'd24;
        rom[352][18] = 8'd3;
        rom[352][19] = 8'd27;
        rom[352][20] = -8'd4;
        rom[352][21] = 8'd5;
        rom[352][22] = -8'd37;
        rom[352][23] = -8'd9;
        rom[352][24] = 8'd3;
        rom[352][25] = -8'd20;
        rom[352][26] = 8'd8;
        rom[352][27] = -8'd26;
        rom[352][28] = 8'd7;
        rom[352][29] = 8'd21;
        rom[352][30] = 8'd24;
        rom[352][31] = -8'd15;
        rom[352][32] = 8'd36;
        rom[352][33] = -8'd11;
        rom[352][34] = -8'd17;
        rom[352][35] = 8'd4;
        rom[352][36] = 8'd6;
        rom[352][37] = 8'd1;
        rom[352][38] = -8'd16;
        rom[352][39] = -8'd33;
        rom[352][40] = 8'd23;
        rom[352][41] = -8'd7;
        rom[352][42] = 8'd40;
        rom[352][43] = -8'd5;
        rom[352][44] = -8'd23;
        rom[352][45] = 8'd19;
        rom[352][46] = -8'd8;
        rom[352][47] = -8'd41;
        rom[352][48] = -8'd12;
        rom[352][49] = -8'd18;
        rom[352][50] = 8'd21;
        rom[352][51] = 8'd2;
        rom[352][52] = -8'd2;
        rom[352][53] = -8'd2;
        rom[352][54] = -8'd35;
        rom[352][55] = 8'd12;
        rom[352][56] = -8'd10;
        rom[352][57] = -8'd11;
        rom[352][58] = 8'd1;
        rom[352][59] = 8'd15;
        rom[352][60] = 8'd63;
        rom[352][61] = -8'd1;
        rom[352][62] = 8'd11;
        rom[352][63] = -8'd5;
        rom[353][0] = -8'd20;
        rom[353][1] = -8'd19;
        rom[353][2] = -8'd8;
        rom[353][3] = -8'd21;
        rom[353][4] = -8'd44;
        rom[353][5] = 8'd1;
        rom[353][6] = 8'd15;
        rom[353][7] = 8'd6;
        rom[353][8] = -8'd11;
        rom[353][9] = -8'd46;
        rom[353][10] = -8'd4;
        rom[353][11] = 8'd2;
        rom[353][12] = 8'd11;
        rom[353][13] = 8'd2;
        rom[353][14] = 8'd30;
        rom[353][15] = 8'd27;
        rom[353][16] = 8'd31;
        rom[353][17] = 8'd18;
        rom[353][18] = 8'd20;
        rom[353][19] = -8'd1;
        rom[353][20] = -8'd6;
        rom[353][21] = 8'd24;
        rom[353][22] = 8'd9;
        rom[353][23] = -8'd14;
        rom[353][24] = 8'd23;
        rom[353][25] = 8'd33;
        rom[353][26] = -8'd1;
        rom[353][27] = 8'd9;
        rom[353][28] = -8'd4;
        rom[353][29] = 8'd28;
        rom[353][30] = 8'd15;
        rom[353][31] = 8'd2;
        rom[353][32] = 8'd0;
        rom[353][33] = 8'd21;
        rom[353][34] = -8'd18;
        rom[353][35] = 8'd32;
        rom[353][36] = -8'd3;
        rom[353][37] = 8'd7;
        rom[353][38] = 8'd13;
        rom[353][39] = -8'd16;
        rom[353][40] = -8'd39;
        rom[353][41] = -8'd32;
        rom[353][42] = -8'd13;
        rom[353][43] = 8'd20;
        rom[353][44] = 8'd30;
        rom[353][45] = 8'd4;
        rom[353][46] = -8'd24;
        rom[353][47] = 8'd19;
        rom[353][48] = -8'd1;
        rom[353][49] = 8'd22;
        rom[353][50] = -8'd4;
        rom[353][51] = 8'd15;
        rom[353][52] = -8'd49;
        rom[353][53] = -8'd31;
        rom[353][54] = -8'd28;
        rom[353][55] = 8'd40;
        rom[353][56] = -8'd1;
        rom[353][57] = -8'd11;
        rom[353][58] = 8'd11;
        rom[353][59] = -8'd38;
        rom[353][60] = -8'd68;
        rom[353][61] = -8'd11;
        rom[353][62] = 8'd52;
        rom[353][63] = -8'd1;
        rom[354][0] = -8'd21;
        rom[354][1] = -8'd6;
        rom[354][2] = -8'd8;
        rom[354][3] = 8'd11;
        rom[354][4] = 8'd2;
        rom[354][5] = 8'd11;
        rom[354][6] = -8'd20;
        rom[354][7] = 8'd11;
        rom[354][8] = 8'd20;
        rom[354][9] = -8'd34;
        rom[354][10] = -8'd13;
        rom[354][11] = -8'd6;
        rom[354][12] = 8'd1;
        rom[354][13] = 8'd23;
        rom[354][14] = -8'd25;
        rom[354][15] = 8'd7;
        rom[354][16] = 8'd12;
        rom[354][17] = -8'd18;
        rom[354][18] = -8'd4;
        rom[354][19] = -8'd5;
        rom[354][20] = -8'd11;
        rom[354][21] = -8'd4;
        rom[354][22] = 8'd29;
        rom[354][23] = 8'd39;
        rom[354][24] = 8'd8;
        rom[354][25] = 8'd25;
        rom[354][26] = -8'd6;
        rom[354][27] = -8'd27;
        rom[354][28] = -8'd38;
        rom[354][29] = -8'd46;
        rom[354][30] = -8'd27;
        rom[354][31] = -8'd22;
        rom[354][32] = -8'd28;
        rom[354][33] = -8'd1;
        rom[354][34] = 8'd16;
        rom[354][35] = -8'd10;
        rom[354][36] = -8'd3;
        rom[354][37] = 8'd13;
        rom[354][38] = -8'd20;
        rom[354][39] = 8'd18;
        rom[354][40] = -8'd22;
        rom[354][41] = 8'd4;
        rom[354][42] = -8'd17;
        rom[354][43] = -8'd17;
        rom[354][44] = -8'd65;
        rom[354][45] = 8'd3;
        rom[354][46] = -8'd6;
        rom[354][47] = -8'd13;
        rom[354][48] = -8'd32;
        rom[354][49] = 8'd23;
        rom[354][50] = 8'd0;
        rom[354][51] = 8'd31;
        rom[354][52] = 8'd2;
        rom[354][53] = -8'd7;
        rom[354][54] = 8'd18;
        rom[354][55] = 8'd3;
        rom[354][56] = 8'd14;
        rom[354][57] = -8'd14;
        rom[354][58] = 8'd1;
        rom[354][59] = -8'd12;
        rom[354][60] = -8'd31;
        rom[354][61] = -8'd19;
        rom[354][62] = 8'd19;
        rom[354][63] = -8'd19;
        rom[355][0] = -8'd59;
        rom[355][1] = 8'd20;
        rom[355][2] = 8'd17;
        rom[355][3] = 8'd48;
        rom[355][4] = -8'd7;
        rom[355][5] = -8'd5;
        rom[355][6] = -8'd15;
        rom[355][7] = -8'd28;
        rom[355][8] = -8'd4;
        rom[355][9] = -8'd67;
        rom[355][10] = 8'd20;
        rom[355][11] = 8'd16;
        rom[355][12] = 8'd44;
        rom[355][13] = -8'd4;
        rom[355][14] = 8'd1;
        rom[355][15] = 8'd11;
        rom[355][16] = 8'd32;
        rom[355][17] = 8'd28;
        rom[355][18] = -8'd17;
        rom[355][19] = -8'd11;
        rom[355][20] = 8'd0;
        rom[355][21] = -8'd18;
        rom[355][22] = -8'd20;
        rom[355][23] = -8'd23;
        rom[355][24] = 8'd19;
        rom[355][25] = -8'd50;
        rom[355][26] = -8'd37;
        rom[355][27] = -8'd8;
        rom[355][28] = 8'd4;
        rom[355][29] = -8'd16;
        rom[355][30] = 8'd31;
        rom[355][31] = -8'd19;
        rom[355][32] = -8'd33;
        rom[355][33] = -8'd13;
        rom[355][34] = 8'd11;
        rom[355][35] = -8'd11;
        rom[355][36] = -8'd13;
        rom[355][37] = 8'd32;
        rom[355][38] = -8'd56;
        rom[355][39] = -8'd7;
        rom[355][40] = -8'd6;
        rom[355][41] = -8'd26;
        rom[355][42] = 8'd8;
        rom[355][43] = 8'd9;
        rom[355][44] = 8'd23;
        rom[355][45] = 8'd5;
        rom[355][46] = 8'd2;
        rom[355][47] = -8'd11;
        rom[355][48] = -8'd1;
        rom[355][49] = 8'd18;
        rom[355][50] = 8'd18;
        rom[355][51] = 8'd10;
        rom[355][52] = -8'd7;
        rom[355][53] = -8'd51;
        rom[355][54] = -8'd30;
        rom[355][55] = -8'd76;
        rom[355][56] = -8'd7;
        rom[355][57] = -8'd16;
        rom[355][58] = 8'd19;
        rom[355][59] = -8'd15;
        rom[355][60] = -8'd76;
        rom[355][61] = -8'd38;
        rom[355][62] = -8'd20;
        rom[355][63] = -8'd15;
        rom[356][0] = -8'd26;
        rom[356][1] = -8'd10;
        rom[356][2] = 8'd13;
        rom[356][3] = 8'd14;
        rom[356][4] = -8'd10;
        rom[356][5] = -8'd10;
        rom[356][6] = -8'd30;
        rom[356][7] = -8'd5;
        rom[356][8] = 8'd4;
        rom[356][9] = -8'd27;
        rom[356][10] = -8'd2;
        rom[356][11] = -8'd1;
        rom[356][12] = 8'd9;
        rom[356][13] = -8'd57;
        rom[356][14] = -8'd5;
        rom[356][15] = -8'd34;
        rom[356][16] = -8'd6;
        rom[356][17] = 8'd22;
        rom[356][18] = 8'd0;
        rom[356][19] = 8'd16;
        rom[356][20] = -8'd2;
        rom[356][21] = -8'd2;
        rom[356][22] = -8'd3;
        rom[356][23] = -8'd33;
        rom[356][24] = -8'd11;
        rom[356][25] = -8'd4;
        rom[356][26] = 8'd22;
        rom[356][27] = 8'd14;
        rom[356][28] = 8'd41;
        rom[356][29] = 8'd2;
        rom[356][30] = -8'd28;
        rom[356][31] = 8'd7;
        rom[356][32] = -8'd31;
        rom[356][33] = -8'd5;
        rom[356][34] = -8'd38;
        rom[356][35] = -8'd52;
        rom[356][36] = -8'd7;
        rom[356][37] = 8'd0;
        rom[356][38] = -8'd12;
        rom[356][39] = -8'd7;
        rom[356][40] = 8'd13;
        rom[356][41] = -8'd6;
        rom[356][42] = -8'd37;
        rom[356][43] = 8'd10;
        rom[356][44] = 8'd17;
        rom[356][45] = -8'd26;
        rom[356][46] = -8'd85;
        rom[356][47] = 8'd1;
        rom[356][48] = -8'd19;
        rom[356][49] = -8'd30;
        rom[356][50] = -8'd4;
        rom[356][51] = -8'd8;
        rom[356][52] = -8'd95;
        rom[356][53] = -8'd11;
        rom[356][54] = -8'd38;
        rom[356][55] = -8'd10;
        rom[356][56] = -8'd5;
        rom[356][57] = 8'd13;
        rom[356][58] = -8'd26;
        rom[356][59] = -8'd34;
        rom[356][60] = -8'd90;
        rom[356][61] = -8'd22;
        rom[356][62] = -8'd16;
        rom[356][63] = -8'd28;
        rom[357][0] = -8'd10;
        rom[357][1] = -8'd69;
        rom[357][2] = 8'd6;
        rom[357][3] = -8'd6;
        rom[357][4] = -8'd50;
        rom[357][5] = 8'd20;
        rom[357][6] = -8'd42;
        rom[357][7] = 8'd1;
        rom[357][8] = -8'd3;
        rom[357][9] = 8'd10;
        rom[357][10] = -8'd15;
        rom[357][11] = 8'd6;
        rom[357][12] = 8'd2;
        rom[357][13] = 8'd15;
        rom[357][14] = -8'd16;
        rom[357][15] = 8'd3;
        rom[357][16] = -8'd76;
        rom[357][17] = 8'd30;
        rom[357][18] = 8'd4;
        rom[357][19] = -8'd65;
        rom[357][20] = -8'd12;
        rom[357][21] = 8'd14;
        rom[357][22] = -8'd15;
        rom[357][23] = 8'd12;
        rom[357][24] = -8'd32;
        rom[357][25] = 8'd21;
        rom[357][26] = -8'd3;
        rom[357][27] = -8'd74;
        rom[357][28] = 8'd8;
        rom[357][29] = 8'd5;
        rom[357][30] = 8'd13;
        rom[357][31] = 8'd15;
        rom[357][32] = -8'd16;
        rom[357][33] = 8'd6;
        rom[357][34] = -8'd10;
        rom[357][35] = -8'd27;
        rom[357][36] = -8'd10;
        rom[357][37] = -8'd22;
        rom[357][38] = -8'd15;
        rom[357][39] = 8'd19;
        rom[357][40] = 8'd10;
        rom[357][41] = -8'd36;
        rom[357][42] = 8'd41;
        rom[357][43] = 8'd11;
        rom[357][44] = 8'd22;
        rom[357][45] = -8'd30;
        rom[357][46] = 8'd27;
        rom[357][47] = 8'd12;
        rom[357][48] = -8'd14;
        rom[357][49] = -8'd20;
        rom[357][50] = -8'd24;
        rom[357][51] = -8'd49;
        rom[357][52] = 8'd25;
        rom[357][53] = 8'd7;
        rom[357][54] = -8'd16;
        rom[357][55] = 8'd14;
        rom[357][56] = -8'd106;
        rom[357][57] = 8'd13;
        rom[357][58] = -8'd43;
        rom[357][59] = 8'd50;
        rom[357][60] = -8'd21;
        rom[357][61] = 8'd11;
        rom[357][62] = 8'd4;
        rom[357][63] = -8'd61;
        rom[358][0] = -8'd20;
        rom[358][1] = -8'd47;
        rom[358][2] = -8'd12;
        rom[358][3] = -8'd49;
        rom[358][4] = -8'd28;
        rom[358][5] = 8'd19;
        rom[358][6] = 8'd4;
        rom[358][7] = 8'd36;
        rom[358][8] = 8'd60;
        rom[358][9] = 8'd26;
        rom[358][10] = -8'd46;
        rom[358][11] = 8'd24;
        rom[358][12] = -8'd6;
        rom[358][13] = -8'd12;
        rom[358][14] = -8'd29;
        rom[358][15] = 8'd2;
        rom[358][16] = 8'd23;
        rom[358][17] = -8'd15;
        rom[358][18] = 8'd7;
        rom[358][19] = -8'd30;
        rom[358][20] = -8'd2;
        rom[358][21] = -8'd31;
        rom[358][22] = -8'd51;
        rom[358][23] = -8'd1;
        rom[358][24] = -8'd32;
        rom[358][25] = 8'd21;
        rom[358][26] = 8'd11;
        rom[358][27] = -8'd59;
        rom[358][28] = 8'd54;
        rom[358][29] = -8'd3;
        rom[358][30] = 8'd43;
        rom[358][31] = 8'd18;
        rom[358][32] = 8'd3;
        rom[358][33] = 8'd30;
        rom[358][34] = -8'd24;
        rom[358][35] = 8'd15;
        rom[358][36] = 8'd46;
        rom[358][37] = 8'd9;
        rom[358][38] = -8'd30;
        rom[358][39] = -8'd16;
        rom[358][40] = 8'd6;
        rom[358][41] = 8'd1;
        rom[358][42] = -8'd59;
        rom[358][43] = 8'd56;
        rom[358][44] = 8'd17;
        rom[358][45] = -8'd4;
        rom[358][46] = 8'd2;
        rom[358][47] = 8'd29;
        rom[358][48] = -8'd15;
        rom[358][49] = -8'd10;
        rom[358][50] = 8'd2;
        rom[358][51] = -8'd42;
        rom[358][52] = 8'd34;
        rom[358][53] = -8'd12;
        rom[358][54] = 8'd2;
        rom[358][55] = -8'd12;
        rom[358][56] = -8'd53;
        rom[358][57] = 8'd11;
        rom[358][58] = -8'd38;
        rom[358][59] = 8'd61;
        rom[358][60] = -8'd5;
        rom[358][61] = 8'd7;
        rom[358][62] = 8'd6;
        rom[358][63] = -8'd3;
        rom[359][0] = 8'd19;
        rom[359][1] = -8'd17;
        rom[359][2] = 8'd18;
        rom[359][3] = -8'd9;
        rom[359][4] = -8'd35;
        rom[359][5] = 8'd17;
        rom[359][6] = 8'd22;
        rom[359][7] = -8'd6;
        rom[359][8] = 8'd34;
        rom[359][9] = 8'd29;
        rom[359][10] = -8'd24;
        rom[359][11] = 8'd36;
        rom[359][12] = -8'd10;
        rom[359][13] = 8'd9;
        rom[359][14] = 8'd39;
        rom[359][15] = 8'd24;
        rom[359][16] = 8'd5;
        rom[359][17] = -8'd29;
        rom[359][18] = 8'd15;
        rom[359][19] = -8'd22;
        rom[359][20] = 8'd0;
        rom[359][21] = -8'd29;
        rom[359][22] = -8'd29;
        rom[359][23] = 8'd41;
        rom[359][24] = -8'd5;
        rom[359][25] = -8'd29;
        rom[359][26] = -8'd5;
        rom[359][27] = 8'd2;
        rom[359][28] = 8'd11;
        rom[359][29] = 8'd45;
        rom[359][30] = 8'd2;
        rom[359][31] = 8'd35;
        rom[359][32] = -8'd28;
        rom[359][33] = 8'd14;
        rom[359][34] = -8'd33;
        rom[359][35] = -8'd10;
        rom[359][36] = -8'd10;
        rom[359][37] = -8'd14;
        rom[359][38] = -8'd2;
        rom[359][39] = 8'd16;
        rom[359][40] = -8'd4;
        rom[359][41] = -8'd59;
        rom[359][42] = 8'd7;
        rom[359][43] = -8'd8;
        rom[359][44] = -8'd34;
        rom[359][45] = -8'd15;
        rom[359][46] = -8'd13;
        rom[359][47] = -8'd57;
        rom[359][48] = 8'd9;
        rom[359][49] = 8'd30;
        rom[359][50] = 8'd42;
        rom[359][51] = 8'd16;
        rom[359][52] = -8'd7;
        rom[359][53] = 8'd12;
        rom[359][54] = -8'd18;
        rom[359][55] = -8'd43;
        rom[359][56] = -8'd2;
        rom[359][57] = 8'd14;
        rom[359][58] = -8'd24;
        rom[359][59] = 8'd39;
        rom[359][60] = 8'd17;
        rom[359][61] = -8'd24;
        rom[359][62] = 8'd3;
        rom[359][63] = 8'd7;
        rom[360][0] = -8'd24;
        rom[360][1] = 8'd7;
        rom[360][2] = -8'd34;
        rom[360][3] = 8'd8;
        rom[360][4] = 8'd13;
        rom[360][5] = -8'd10;
        rom[360][6] = 8'd29;
        rom[360][7] = -8'd4;
        rom[360][8] = -8'd10;
        rom[360][9] = -8'd31;
        rom[360][10] = 8'd44;
        rom[360][11] = -8'd28;
        rom[360][12] = -8'd40;
        rom[360][13] = 8'd44;
        rom[360][14] = -8'd3;
        rom[360][15] = -8'd70;
        rom[360][16] = -8'd30;
        rom[360][17] = 8'd5;
        rom[360][18] = -8'd5;
        rom[360][19] = -8'd3;
        rom[360][20] = 8'd6;
        rom[360][21] = 8'd25;
        rom[360][22] = 8'd14;
        rom[360][23] = -8'd9;
        rom[360][24] = -8'd39;
        rom[360][25] = 8'd9;
        rom[360][26] = 8'd1;
        rom[360][27] = -8'd19;
        rom[360][28] = 8'd26;
        rom[360][29] = -8'd38;
        rom[360][30] = 8'd10;
        rom[360][31] = -8'd17;
        rom[360][32] = 8'd15;
        rom[360][33] = 8'd12;
        rom[360][34] = -8'd14;
        rom[360][35] = -8'd19;
        rom[360][36] = 8'd11;
        rom[360][37] = -8'd9;
        rom[360][38] = 8'd21;
        rom[360][39] = 8'd36;
        rom[360][40] = -8'd8;
        rom[360][41] = 8'd7;
        rom[360][42] = -8'd42;
        rom[360][43] = 8'd13;
        rom[360][44] = 8'd21;
        rom[360][45] = -8'd18;
        rom[360][46] = -8'd31;
        rom[360][47] = -8'd17;
        rom[360][48] = -8'd5;
        rom[360][49] = 8'd1;
        rom[360][50] = 8'd19;
        rom[360][51] = -8'd34;
        rom[360][52] = -8'd18;
        rom[360][53] = -8'd13;
        rom[360][54] = -8'd11;
        rom[360][55] = -8'd20;
        rom[360][56] = 8'd60;
        rom[360][57] = 8'd38;
        rom[360][58] = 8'd15;
        rom[360][59] = -8'd71;
        rom[360][60] = 8'd26;
        rom[360][61] = -8'd31;
        rom[360][62] = -8'd19;
        rom[360][63] = 8'd27;
        rom[361][0] = 8'd20;
        rom[361][1] = 8'd8;
        rom[361][2] = 8'd7;
        rom[361][3] = -8'd2;
        rom[361][4] = -8'd2;
        rom[361][5] = -8'd10;
        rom[361][6] = 8'd18;
        rom[361][7] = -8'd20;
        rom[361][8] = 8'd9;
        rom[361][9] = 8'd8;
        rom[361][10] = -8'd30;
        rom[361][11] = -8'd12;
        rom[361][12] = -8'd48;
        rom[361][13] = -8'd33;
        rom[361][14] = -8'd25;
        rom[361][15] = 8'd17;
        rom[361][16] = -8'd37;
        rom[361][17] = 8'd6;
        rom[361][18] = 8'd10;
        rom[361][19] = -8'd3;
        rom[361][20] = -8'd2;
        rom[361][21] = 8'd29;
        rom[361][22] = 8'd11;
        rom[361][23] = -8'd25;
        rom[361][24] = -8'd47;
        rom[361][25] = 8'd34;
        rom[361][26] = 8'd18;
        rom[361][27] = -8'd33;
        rom[361][28] = -8'd1;
        rom[361][29] = -8'd21;
        rom[361][30] = 8'd24;
        rom[361][31] = 8'd17;
        rom[361][32] = 8'd7;
        rom[361][33] = 8'd20;
        rom[361][34] = 8'd5;
        rom[361][35] = 8'd10;
        rom[361][36] = 8'd1;
        rom[361][37] = -8'd26;
        rom[361][38] = 8'd10;
        rom[361][39] = -8'd49;
        rom[361][40] = 8'd2;
        rom[361][41] = 8'd44;
        rom[361][42] = -8'd23;
        rom[361][43] = 8'd29;
        rom[361][44] = 8'd14;
        rom[361][45] = -8'd52;
        rom[361][46] = -8'd17;
        rom[361][47] = -8'd12;
        rom[361][48] = -8'd17;
        rom[361][49] = 8'd0;
        rom[361][50] = -8'd16;
        rom[361][51] = 8'd16;
        rom[361][52] = -8'd1;
        rom[361][53] = 8'd27;
        rom[361][54] = 8'd35;
        rom[361][55] = 8'd30;
        rom[361][56] = 8'd6;
        rom[361][57] = -8'd30;
        rom[361][58] = -8'd4;
        rom[361][59] = -8'd31;
        rom[361][60] = 8'd7;
        rom[361][61] = -8'd66;
        rom[361][62] = -8'd14;
        rom[361][63] = -8'd20;
        rom[362][0] = -8'd40;
        rom[362][1] = 8'd15;
        rom[362][2] = 8'd3;
        rom[362][3] = -8'd43;
        rom[362][4] = -8'd8;
        rom[362][5] = -8'd15;
        rom[362][6] = -8'd1;
        rom[362][7] = 8'd19;
        rom[362][8] = 8'd5;
        rom[362][9] = 8'd5;
        rom[362][10] = -8'd19;
        rom[362][11] = 8'd8;
        rom[362][12] = 8'd8;
        rom[362][13] = 8'd32;
        rom[362][14] = -8'd28;
        rom[362][15] = -8'd47;
        rom[362][16] = 8'd35;
        rom[362][17] = -8'd59;
        rom[362][18] = -8'd8;
        rom[362][19] = -8'd14;
        rom[362][20] = 8'd6;
        rom[362][21] = 8'd13;
        rom[362][22] = -8'd10;
        rom[362][23] = 8'd16;
        rom[362][24] = -8'd45;
        rom[362][25] = -8'd11;
        rom[362][26] = -8'd49;
        rom[362][27] = -8'd92;
        rom[362][28] = 8'd3;
        rom[362][29] = 8'd15;
        rom[362][30] = -8'd10;
        rom[362][31] = 8'd34;
        rom[362][32] = 8'd27;
        rom[362][33] = 8'd23;
        rom[362][34] = -8'd51;
        rom[362][35] = -8'd22;
        rom[362][36] = -8'd31;
        rom[362][37] = 8'd3;
        rom[362][38] = -8'd25;
        rom[362][39] = 8'd5;
        rom[362][40] = -8'd9;
        rom[362][41] = 8'd5;
        rom[362][42] = -8'd9;
        rom[362][43] = 8'd1;
        rom[362][44] = -8'd38;
        rom[362][45] = 8'd5;
        rom[362][46] = 8'd27;
        rom[362][47] = 8'd20;
        rom[362][48] = -8'd15;
        rom[362][49] = -8'd1;
        rom[362][50] = 8'd6;
        rom[362][51] = -8'd37;
        rom[362][52] = -8'd14;
        rom[362][53] = -8'd21;
        rom[362][54] = 8'd4;
        rom[362][55] = 8'd22;
        rom[362][56] = -8'd20;
        rom[362][57] = -8'd18;
        rom[362][58] = -8'd7;
        rom[362][59] = -8'd13;
        rom[362][60] = -8'd16;
        rom[362][61] = 8'd28;
        rom[362][62] = 8'd22;
        rom[362][63] = 8'd11;
        rom[363][0] = -8'd32;
        rom[363][1] = -8'd12;
        rom[363][2] = -8'd37;
        rom[363][3] = 8'd3;
        rom[363][4] = -8'd28;
        rom[363][5] = -8'd33;
        rom[363][6] = -8'd5;
        rom[363][7] = -8'd5;
        rom[363][8] = -8'd22;
        rom[363][9] = 8'd17;
        rom[363][10] = -8'd60;
        rom[363][11] = 8'd6;
        rom[363][12] = -8'd56;
        rom[363][13] = 8'd7;
        rom[363][14] = -8'd52;
        rom[363][15] = -8'd49;
        rom[363][16] = -8'd45;
        rom[363][17] = -8'd49;
        rom[363][18] = -8'd18;
        rom[363][19] = 8'd10;
        rom[363][20] = -8'd7;
        rom[363][21] = -8'd6;
        rom[363][22] = 8'd5;
        rom[363][23] = -8'd21;
        rom[363][24] = -8'd6;
        rom[363][25] = -8'd23;
        rom[363][26] = 8'd0;
        rom[363][27] = -8'd65;
        rom[363][28] = -8'd20;
        rom[363][29] = -8'd24;
        rom[363][30] = -8'd7;
        rom[363][31] = 8'd13;
        rom[363][32] = -8'd13;
        rom[363][33] = -8'd16;
        rom[363][34] = -8'd27;
        rom[363][35] = -8'd10;
        rom[363][36] = -8'd12;
        rom[363][37] = -8'd16;
        rom[363][38] = 8'd42;
        rom[363][39] = 8'd1;
        rom[363][40] = -8'd20;
        rom[363][41] = 8'd5;
        rom[363][42] = -8'd26;
        rom[363][43] = -8'd9;
        rom[363][44] = 8'd9;
        rom[363][45] = 8'd26;
        rom[363][46] = 8'd10;
        rom[363][47] = 8'd11;
        rom[363][48] = -8'd34;
        rom[363][49] = -8'd46;
        rom[363][50] = -8'd25;
        rom[363][51] = 8'd44;
        rom[363][52] = -8'd5;
        rom[363][53] = -8'd17;
        rom[363][54] = 8'd37;
        rom[363][55] = -8'd52;
        rom[363][56] = -8'd37;
        rom[363][57] = -8'd45;
        rom[363][58] = -8'd2;
        rom[363][59] = 8'd3;
        rom[363][60] = -8'd14;
        rom[363][61] = -8'd5;
        rom[363][62] = -8'd47;
        rom[363][63] = -8'd6;
        rom[364][0] = -8'd14;
        rom[364][1] = -8'd55;
        rom[364][2] = 8'd8;
        rom[364][3] = -8'd26;
        rom[364][4] = -8'd6;
        rom[364][5] = 8'd20;
        rom[364][6] = -8'd11;
        rom[364][7] = -8'd27;
        rom[364][8] = -8'd10;
        rom[364][9] = -8'd16;
        rom[364][10] = -8'd50;
        rom[364][11] = -8'd48;
        rom[364][12] = 8'd7;
        rom[364][13] = -8'd13;
        rom[364][14] = -8'd32;
        rom[364][15] = 8'd26;
        rom[364][16] = -8'd49;
        rom[364][17] = 8'd13;
        rom[364][18] = 8'd17;
        rom[364][19] = 8'd0;
        rom[364][20] = -8'd9;
        rom[364][21] = -8'd3;
        rom[364][22] = -8'd55;
        rom[364][23] = -8'd12;
        rom[364][24] = -8'd60;
        rom[364][25] = -8'd13;
        rom[364][26] = -8'd48;
        rom[364][27] = -8'd63;
        rom[364][28] = -8'd31;
        rom[364][29] = -8'd23;
        rom[364][30] = -8'd12;
        rom[364][31] = 8'd5;
        rom[364][32] = -8'd45;
        rom[364][33] = 8'd0;
        rom[364][34] = -8'd18;
        rom[364][35] = -8'd15;
        rom[364][36] = 8'd23;
        rom[364][37] = -8'd8;
        rom[364][38] = -8'd55;
        rom[364][39] = 8'd31;
        rom[364][40] = -8'd44;
        rom[364][41] = -8'd32;
        rom[364][42] = -8'd41;
        rom[364][43] = -8'd28;
        rom[364][44] = 8'd26;
        rom[364][45] = 8'd4;
        rom[364][46] = 8'd8;
        rom[364][47] = -8'd10;
        rom[364][48] = -8'd3;
        rom[364][49] = 8'd7;
        rom[364][50] = -8'd13;
        rom[364][51] = -8'd38;
        rom[364][52] = -8'd30;
        rom[364][53] = 8'd37;
        rom[364][54] = 8'd19;
        rom[364][55] = -8'd12;
        rom[364][56] = -8'd76;
        rom[364][57] = -8'd7;
        rom[364][58] = -8'd17;
        rom[364][59] = -8'd35;
        rom[364][60] = -8'd1;
        rom[364][61] = -8'd6;
        rom[364][62] = -8'd30;
        rom[364][63] = 8'd19;
        rom[365][0] = 8'd15;
        rom[365][1] = -8'd49;
        rom[365][2] = 8'd22;
        rom[365][3] = 8'd13;
        rom[365][4] = 8'd4;
        rom[365][5] = -8'd4;
        rom[365][6] = -8'd21;
        rom[365][7] = 8'd8;
        rom[365][8] = -8'd6;
        rom[365][9] = -8'd21;
        rom[365][10] = 8'd60;
        rom[365][11] = 8'd47;
        rom[365][12] = 8'd56;
        rom[365][13] = 8'd31;
        rom[365][14] = -8'd6;
        rom[365][15] = -8'd11;
        rom[365][16] = 8'd2;
        rom[365][17] = 8'd2;
        rom[365][18] = -8'd36;
        rom[365][19] = 8'd13;
        rom[365][20] = -8'd8;
        rom[365][21] = 8'd22;
        rom[365][22] = -8'd28;
        rom[365][23] = -8'd27;
        rom[365][24] = 8'd23;
        rom[365][25] = -8'd40;
        rom[365][26] = 8'd23;
        rom[365][27] = 8'd64;
        rom[365][28] = 8'd12;
        rom[365][29] = 8'd4;
        rom[365][30] = -8'd1;
        rom[365][31] = 8'd4;
        rom[365][32] = 8'd7;
        rom[365][33] = -8'd50;
        rom[365][34] = -8'd5;
        rom[365][35] = -8'd38;
        rom[365][36] = -8'd17;
        rom[365][37] = -8'd19;
        rom[365][38] = 8'd21;
        rom[365][39] = -8'd18;
        rom[365][40] = -8'd6;
        rom[365][41] = -8'd39;
        rom[365][42] = 8'd36;
        rom[365][43] = -8'd9;
        rom[365][44] = 8'd12;
        rom[365][45] = -8'd36;
        rom[365][46] = 8'd10;
        rom[365][47] = -8'd41;
        rom[365][48] = -8'd6;
        rom[365][49] = -8'd21;
        rom[365][50] = 8'd19;
        rom[365][51] = -8'd5;
        rom[365][52] = -8'd59;
        rom[365][53] = 8'd16;
        rom[365][54] = -8'd8;
        rom[365][55] = -8'd10;
        rom[365][56] = -8'd5;
        rom[365][57] = -8'd47;
        rom[365][58] = -8'd88;
        rom[365][59] = 8'd26;
        rom[365][60] = 8'd30;
        rom[365][61] = 8'd34;
        rom[365][62] = -8'd4;
        rom[365][63] = -8'd26;
        rom[366][0] = -8'd13;
        rom[366][1] = -8'd19;
        rom[366][2] = 8'd2;
        rom[366][3] = 8'd30;
        rom[366][4] = 8'd16;
        rom[366][5] = 8'd10;
        rom[366][6] = 8'd11;
        rom[366][7] = 8'd32;
        rom[366][8] = -8'd3;
        rom[366][9] = -8'd20;
        rom[366][10] = -8'd25;
        rom[366][11] = 8'd8;
        rom[366][12] = -8'd12;
        rom[366][13] = 8'd4;
        rom[366][14] = 8'd8;
        rom[366][15] = 8'd15;
        rom[366][16] = -8'd17;
        rom[366][17] = 8'd9;
        rom[366][18] = 8'd18;
        rom[366][19] = 8'd13;
        rom[366][20] = -8'd7;
        rom[366][21] = -8'd10;
        rom[366][22] = 8'd35;
        rom[366][23] = 8'd7;
        rom[366][24] = -8'd52;
        rom[366][25] = 8'd4;
        rom[366][26] = -8'd2;
        rom[366][27] = -8'd17;
        rom[366][28] = 8'd12;
        rom[366][29] = -8'd1;
        rom[366][30] = -8'd4;
        rom[366][31] = 8'd15;
        rom[366][32] = 8'd9;
        rom[366][33] = 8'd35;
        rom[366][34] = 8'd18;
        rom[366][35] = 8'd23;
        rom[366][36] = 8'd41;
        rom[366][37] = -8'd29;
        rom[366][38] = -8'd48;
        rom[366][39] = -8'd15;
        rom[366][40] = -8'd7;
        rom[366][41] = 8'd3;
        rom[366][42] = 8'd11;
        rom[366][43] = 8'd1;
        rom[366][44] = 8'd39;
        rom[366][45] = 8'd2;
        rom[366][46] = 8'd7;
        rom[366][47] = 8'd4;
        rom[366][48] = -8'd7;
        rom[366][49] = 8'd41;
        rom[366][50] = -8'd23;
        rom[366][51] = 8'd0;
        rom[366][52] = 8'd19;
        rom[366][53] = -8'd18;
        rom[366][54] = 8'd8;
        rom[366][55] = 8'd35;
        rom[366][56] = 8'd11;
        rom[366][57] = 8'd1;
        rom[366][58] = -8'd6;
        rom[366][59] = -8'd39;
        rom[366][60] = -8'd33;
        rom[366][61] = -8'd23;
        rom[366][62] = -8'd58;
        rom[366][63] = -8'd56;
        rom[367][0] = -8'd45;
        rom[367][1] = -8'd3;
        rom[367][2] = -8'd99;
        rom[367][3] = 8'd7;
        rom[367][4] = -8'd3;
        rom[367][5] = 8'd5;
        rom[367][6] = 8'd15;
        rom[367][7] = -8'd26;
        rom[367][8] = -8'd53;
        rom[367][9] = -8'd69;
        rom[367][10] = 8'd24;
        rom[367][11] = 8'd37;
        rom[367][12] = 8'd9;
        rom[367][13] = 8'd5;
        rom[367][14] = 8'd13;
        rom[367][15] = -8'd34;
        rom[367][16] = 8'd15;
        rom[367][17] = 8'd44;
        rom[367][18] = -8'd30;
        rom[367][19] = 8'd52;
        rom[367][20] = 8'd2;
        rom[367][21] = -8'd15;
        rom[367][22] = 8'd9;
        rom[367][23] = -8'd5;
        rom[367][24] = -8'd16;
        rom[367][25] = 8'd17;
        rom[367][26] = -8'd24;
        rom[367][27] = 8'd55;
        rom[367][28] = -8'd39;
        rom[367][29] = -8'd2;
        rom[367][30] = 8'd18;
        rom[367][31] = 8'd52;
        rom[367][32] = 8'd16;
        rom[367][33] = -8'd4;
        rom[367][34] = -8'd13;
        rom[367][35] = 8'd37;
        rom[367][36] = -8'd8;
        rom[367][37] = 8'd17;
        rom[367][38] = -8'd13;
        rom[367][39] = 8'd10;
        rom[367][40] = -8'd22;
        rom[367][41] = 8'd30;
        rom[367][42] = -8'd13;
        rom[367][43] = 8'd34;
        rom[367][44] = 8'd48;
        rom[367][45] = 8'd3;
        rom[367][46] = -8'd60;
        rom[367][47] = -8'd1;
        rom[367][48] = -8'd15;
        rom[367][49] = 8'd2;
        rom[367][50] = 8'd11;
        rom[367][51] = -8'd25;
        rom[367][52] = -8'd21;
        rom[367][53] = -8'd5;
        rom[367][54] = 8'd27;
        rom[367][55] = -8'd11;
        rom[367][56] = -8'd10;
        rom[367][57] = -8'd38;
        rom[367][58] = -8'd17;
        rom[367][59] = -8'd44;
        rom[367][60] = 8'd1;
        rom[367][61] = -8'd25;
        rom[367][62] = -8'd18;
        rom[367][63] = 8'd16;
        rom[368][0] = -8'd12;
        rom[368][1] = 8'd54;
        rom[368][2] = -8'd10;
        rom[368][3] = -8'd16;
        rom[368][4] = -8'd11;
        rom[368][5] = -8'd1;
        rom[368][6] = -8'd78;
        rom[368][7] = -8'd21;
        rom[368][8] = -8'd32;
        rom[368][9] = 8'd11;
        rom[368][10] = -8'd24;
        rom[368][11] = -8'd17;
        rom[368][12] = 8'd26;
        rom[368][13] = -8'd27;
        rom[368][14] = -8'd4;
        rom[368][15] = 8'd30;
        rom[368][16] = 8'd21;
        rom[368][17] = 8'd6;
        rom[368][18] = -8'd27;
        rom[368][19] = -8'd6;
        rom[368][20] = -8'd16;
        rom[368][21] = -8'd10;
        rom[368][22] = -8'd29;
        rom[368][23] = -8'd25;
        rom[368][24] = 8'd0;
        rom[368][25] = -8'd31;
        rom[368][26] = -8'd3;
        rom[368][27] = 8'd9;
        rom[368][28] = -8'd43;
        rom[368][29] = -8'd52;
        rom[368][30] = -8'd23;
        rom[368][31] = -8'd8;
        rom[368][32] = 8'd0;
        rom[368][33] = 8'd34;
        rom[368][34] = -8'd13;
        rom[368][35] = 8'd35;
        rom[368][36] = -8'd34;
        rom[368][37] = 8'd6;
        rom[368][38] = -8'd52;
        rom[368][39] = -8'd17;
        rom[368][40] = 8'd12;
        rom[368][41] = -8'd11;
        rom[368][42] = -8'd7;
        rom[368][43] = 8'd15;
        rom[368][44] = 8'd30;
        rom[368][45] = 8'd28;
        rom[368][46] = 8'd34;
        rom[368][47] = 8'd40;
        rom[368][48] = -8'd60;
        rom[368][49] = 8'd4;
        rom[368][50] = 8'd4;
        rom[368][51] = -8'd28;
        rom[368][52] = -8'd1;
        rom[368][53] = -8'd36;
        rom[368][54] = -8'd9;
        rom[368][55] = -8'd14;
        rom[368][56] = 8'd18;
        rom[368][57] = -8'd22;
        rom[368][58] = -8'd23;
        rom[368][59] = -8'd22;
        rom[368][60] = -8'd33;
        rom[368][61] = 8'd1;
        rom[368][62] = 8'd6;
        rom[368][63] = -8'd32;
        rom[369][0] = -8'd23;
        rom[369][1] = -8'd35;
        rom[369][2] = -8'd24;
        rom[369][3] = -8'd44;
        rom[369][4] = -8'd13;
        rom[369][5] = 8'd19;
        rom[369][6] = -8'd16;
        rom[369][7] = -8'd54;
        rom[369][8] = 8'd6;
        rom[369][9] = -8'd10;
        rom[369][10] = -8'd55;
        rom[369][11] = 8'd31;
        rom[369][12] = 8'd14;
        rom[369][13] = 8'd52;
        rom[369][14] = -8'd4;
        rom[369][15] = -8'd24;
        rom[369][16] = -8'd2;
        rom[369][17] = -8'd21;
        rom[369][18] = -8'd1;
        rom[369][19] = -8'd5;
        rom[369][20] = -8'd5;
        rom[369][21] = -8'd17;
        rom[369][22] = -8'd13;
        rom[369][23] = -8'd21;
        rom[369][24] = 8'd39;
        rom[369][25] = -8'd14;
        rom[369][26] = -8'd24;
        rom[369][27] = -8'd27;
        rom[369][28] = 8'd25;
        rom[369][29] = -8'd17;
        rom[369][30] = 8'd43;
        rom[369][31] = 8'd4;
        rom[369][32] = -8'd1;
        rom[369][33] = -8'd24;
        rom[369][34] = -8'd4;
        rom[369][35] = -8'd17;
        rom[369][36] = 8'd33;
        rom[369][37] = -8'd18;
        rom[369][38] = -8'd8;
        rom[369][39] = -8'd49;
        rom[369][40] = -8'd24;
        rom[369][41] = -8'd1;
        rom[369][42] = -8'd40;
        rom[369][43] = 8'd3;
        rom[369][44] = -8'd12;
        rom[369][45] = 8'd7;
        rom[369][46] = -8'd27;
        rom[369][47] = -8'd6;
        rom[369][48] = -8'd23;
        rom[369][49] = 8'd18;
        rom[369][50] = 8'd8;
        rom[369][51] = 8'd42;
        rom[369][52] = -8'd10;
        rom[369][53] = 8'd26;
        rom[369][54] = 8'd37;
        rom[369][55] = 8'd12;
        rom[369][56] = -8'd37;
        rom[369][57] = 8'd8;
        rom[369][58] = -8'd33;
        rom[369][59] = 8'd42;
        rom[369][60] = 8'd38;
        rom[369][61] = -8'd7;
        rom[369][62] = -8'd22;
        rom[369][63] = 8'd14;
        rom[370][0] = -8'd3;
        rom[370][1] = -8'd13;
        rom[370][2] = 8'd15;
        rom[370][3] = -8'd14;
        rom[370][4] = -8'd16;
        rom[370][5] = 8'd9;
        rom[370][6] = 8'd11;
        rom[370][7] = -8'd28;
        rom[370][8] = -8'd10;
        rom[370][9] = -8'd20;
        rom[370][10] = -8'd12;
        rom[370][11] = 8'd18;
        rom[370][12] = 8'd18;
        rom[370][13] = 8'd9;
        rom[370][14] = 8'd6;
        rom[370][15] = -8'd59;
        rom[370][16] = -8'd68;
        rom[370][17] = -8'd26;
        rom[370][18] = -8'd13;
        rom[370][19] = -8'd17;
        rom[370][20] = -8'd8;
        rom[370][21] = 8'd7;
        rom[370][22] = 8'd20;
        rom[370][23] = 8'd33;
        rom[370][24] = 8'd5;
        rom[370][25] = -8'd21;
        rom[370][26] = -8'd34;
        rom[370][27] = 8'd19;
        rom[370][28] = -8'd11;
        rom[370][29] = 8'd14;
        rom[370][30] = -8'd4;
        rom[370][31] = 8'd1;
        rom[370][32] = 8'd39;
        rom[370][33] = -8'd21;
        rom[370][34] = 8'd38;
        rom[370][35] = 8'd24;
        rom[370][36] = -8'd8;
        rom[370][37] = 8'd38;
        rom[370][38] = 8'd3;
        rom[370][39] = 8'd25;
        rom[370][40] = -8'd52;
        rom[370][41] = -8'd3;
        rom[370][42] = -8'd12;
        rom[370][43] = -8'd4;
        rom[370][44] = 8'd6;
        rom[370][45] = 8'd3;
        rom[370][46] = -8'd19;
        rom[370][47] = 8'd18;
        rom[370][48] = 8'd25;
        rom[370][49] = 8'd23;
        rom[370][50] = -8'd8;
        rom[370][51] = -8'd29;
        rom[370][52] = 8'd6;
        rom[370][53] = -8'd44;
        rom[370][54] = -8'd30;
        rom[370][55] = -8'd8;
        rom[370][56] = 8'd16;
        rom[370][57] = 8'd6;
        rom[370][58] = -8'd6;
        rom[370][59] = -8'd42;
        rom[370][60] = -8'd23;
        rom[370][61] = -8'd4;
        rom[370][62] = -8'd17;
        rom[370][63] = 8'd3;
        rom[371][0] = -8'd9;
        rom[371][1] = 8'd7;
        rom[371][2] = 8'd6;
        rom[371][3] = -8'd18;
        rom[371][4] = 8'd10;
        rom[371][5] = -8'd49;
        rom[371][6] = 8'd4;
        rom[371][7] = -8'd30;
        rom[371][8] = 8'd34;
        rom[371][9] = 8'd10;
        rom[371][10] = 8'd24;
        rom[371][11] = 8'd21;
        rom[371][12] = -8'd2;
        rom[371][13] = -8'd37;
        rom[371][14] = 8'd11;
        rom[371][15] = 8'd19;
        rom[371][16] = -8'd11;
        rom[371][17] = 8'd5;
        rom[371][18] = -8'd42;
        rom[371][19] = -8'd6;
        rom[371][20] = 8'd5;
        rom[371][21] = 8'd25;
        rom[371][22] = 8'd9;
        rom[371][23] = -8'd41;
        rom[371][24] = -8'd9;
        rom[371][25] = 8'd2;
        rom[371][26] = -8'd20;
        rom[371][27] = -8'd24;
        rom[371][28] = -8'd30;
        rom[371][29] = 8'd15;
        rom[371][30] = 8'd10;
        rom[371][31] = -8'd15;
        rom[371][32] = -8'd23;
        rom[371][33] = -8'd38;
        rom[371][34] = 8'd17;
        rom[371][35] = -8'd32;
        rom[371][36] = -8'd9;
        rom[371][37] = 8'd46;
        rom[371][38] = -8'd11;
        rom[371][39] = -8'd7;
        rom[371][40] = -8'd39;
        rom[371][41] = -8'd38;
        rom[371][42] = -8'd19;
        rom[371][43] = -8'd37;
        rom[371][44] = 8'd10;
        rom[371][45] = -8'd28;
        rom[371][46] = -8'd8;
        rom[371][47] = -8'd13;
        rom[371][48] = -8'd4;
        rom[371][49] = 8'd9;
        rom[371][50] = -8'd24;
        rom[371][51] = -8'd25;
        rom[371][52] = -8'd25;
        rom[371][53] = 8'd9;
        rom[371][54] = 8'd16;
        rom[371][55] = 8'd30;
        rom[371][56] = -8'd7;
        rom[371][57] = 8'd2;
        rom[371][58] = 8'd5;
        rom[371][59] = -8'd20;
        rom[371][60] = 8'd19;
        rom[371][61] = 8'd40;
        rom[371][62] = 8'd15;
        rom[371][63] = -8'd9;
        rom[372][0] = -8'd24;
        rom[372][1] = -8'd11;
        rom[372][2] = -8'd20;
        rom[372][3] = -8'd3;
        rom[372][4] = 8'd18;
        rom[372][5] = -8'd13;
        rom[372][6] = -8'd97;
        rom[372][7] = -8'd30;
        rom[372][8] = -8'd35;
        rom[372][9] = -8'd43;
        rom[372][10] = -8'd15;
        rom[372][11] = 8'd12;
        rom[372][12] = -8'd68;
        rom[372][13] = -8'd8;
        rom[372][14] = -8'd10;
        rom[372][15] = -8'd60;
        rom[372][16] = -8'd30;
        rom[372][17] = 8'd7;
        rom[372][18] = -8'd6;
        rom[372][19] = -8'd26;
        rom[372][20] = 8'd3;
        rom[372][21] = -8'd43;
        rom[372][22] = -8'd52;
        rom[372][23] = -8'd46;
        rom[372][24] = -8'd24;
        rom[372][25] = -8'd14;
        rom[372][26] = -8'd7;
        rom[372][27] = 8'd19;
        rom[372][28] = -8'd3;
        rom[372][29] = -8'd16;
        rom[372][30] = -8'd20;
        rom[372][31] = -8'd22;
        rom[372][32] = -8'd47;
        rom[372][33] = -8'd2;
        rom[372][34] = -8'd8;
        rom[372][35] = 8'd32;
        rom[372][36] = -8'd31;
        rom[372][37] = -8'd8;
        rom[372][38] = -8'd29;
        rom[372][39] = 8'd33;
        rom[372][40] = 8'd21;
        rom[372][41] = 8'd16;
        rom[372][42] = -8'd32;
        rom[372][43] = -8'd67;
        rom[372][44] = 8'd7;
        rom[372][45] = -8'd2;
        rom[372][46] = -8'd28;
        rom[372][47] = -8'd10;
        rom[372][48] = 8'd5;
        rom[372][49] = 8'd30;
        rom[372][50] = -8'd43;
        rom[372][51] = -8'd6;
        rom[372][52] = -8'd9;
        rom[372][53] = 8'd17;
        rom[372][54] = -8'd52;
        rom[372][55] = 8'd1;
        rom[372][56] = 8'd41;
        rom[372][57] = 8'd3;
        rom[372][58] = -8'd15;
        rom[372][59] = -8'd33;
        rom[372][60] = -8'd9;
        rom[372][61] = -8'd1;
        rom[372][62] = 8'd4;
        rom[372][63] = -8'd15;
        rom[373][0] = -8'd16;
        rom[373][1] = 8'd16;
        rom[373][2] = -8'd57;
        rom[373][3] = -8'd23;
        rom[373][4] = 8'd9;
        rom[373][5] = -8'd46;
        rom[373][6] = 8'd18;
        rom[373][7] = -8'd10;
        rom[373][8] = -8'd12;
        rom[373][9] = 8'd11;
        rom[373][10] = 8'd22;
        rom[373][11] = -8'd6;
        rom[373][12] = 8'd39;
        rom[373][13] = -8'd20;
        rom[373][14] = 8'd35;
        rom[373][15] = -8'd22;
        rom[373][16] = 8'd40;
        rom[373][17] = -8'd43;
        rom[373][18] = 8'd6;
        rom[373][19] = -8'd54;
        rom[373][20] = 8'd2;
        rom[373][21] = 8'd36;
        rom[373][22] = 8'd50;
        rom[373][23] = -8'd24;
        rom[373][24] = -8'd13;
        rom[373][25] = -8'd3;
        rom[373][26] = -8'd21;
        rom[373][27] = -8'd57;
        rom[373][28] = -8'd19;
        rom[373][29] = -8'd29;
        rom[373][30] = -8'd14;
        rom[373][31] = 8'd12;
        rom[373][32] = -8'd14;
        rom[373][33] = -8'd50;
        rom[373][34] = -8'd45;
        rom[373][35] = -8'd11;
        rom[373][36] = -8'd34;
        rom[373][37] = -8'd8;
        rom[373][38] = 8'd9;
        rom[373][39] = 8'd16;
        rom[373][40] = 8'd9;
        rom[373][41] = 8'd14;
        rom[373][42] = -8'd6;
        rom[373][43] = -8'd22;
        rom[373][44] = 8'd6;
        rom[373][45] = 8'd7;
        rom[373][46] = -8'd10;
        rom[373][47] = 8'd18;
        rom[373][48] = -8'd21;
        rom[373][49] = 8'd15;
        rom[373][50] = -8'd31;
        rom[373][51] = -8'd3;
        rom[373][52] = -8'd4;
        rom[373][53] = 8'd13;
        rom[373][54] = 8'd4;
        rom[373][55] = -8'd80;
        rom[373][56] = 8'd8;
        rom[373][57] = 8'd6;
        rom[373][58] = -8'd22;
        rom[373][59] = -8'd36;
        rom[373][60] = 8'd42;
        rom[373][61] = -8'd17;
        rom[373][62] = -8'd29;
        rom[373][63] = -8'd1;
        rom[374][0] = -8'd4;
        rom[374][1] = 8'd8;
        rom[374][2] = -8'd4;
        rom[374][3] = -8'd3;
        rom[374][4] = -8'd9;
        rom[374][5] = 8'd7;
        rom[374][6] = -8'd2;
        rom[374][7] = -8'd11;
        rom[374][8] = 8'd2;
        rom[374][9] = 8'd8;
        rom[374][10] = -8'd4;
        rom[374][11] = -8'd5;
        rom[374][12] = -8'd7;
        rom[374][13] = 8'd7;
        rom[374][14] = 8'd6;
        rom[374][15] = 8'd3;
        rom[374][16] = 8'd0;
        rom[374][17] = 8'd6;
        rom[374][18] = -8'd8;
        rom[374][19] = 8'd7;
        rom[374][20] = 8'd6;
        rom[374][21] = -8'd5;
        rom[374][22] = 8'd3;
        rom[374][23] = 8'd7;
        rom[374][24] = 8'd0;
        rom[374][25] = -8'd10;
        rom[374][26] = -8'd5;
        rom[374][27] = -8'd3;
        rom[374][28] = -8'd4;
        rom[374][29] = -8'd4;
        rom[374][30] = -8'd3;
        rom[374][31] = 8'd4;
        rom[374][32] = -8'd3;
        rom[374][33] = -8'd1;
        rom[374][34] = -8'd1;
        rom[374][35] = 8'd13;
        rom[374][36] = -8'd6;
        rom[374][37] = 8'd6;
        rom[374][38] = -8'd11;
        rom[374][39] = -8'd6;
        rom[374][40] = 8'd2;
        rom[374][41] = -8'd5;
        rom[374][42] = 8'd0;
        rom[374][43] = 8'd0;
        rom[374][44] = 8'd2;
        rom[374][45] = -8'd9;
        rom[374][46] = -8'd2;
        rom[374][47] = -8'd6;
        rom[374][48] = -8'd3;
        rom[374][49] = 8'd4;
        rom[374][50] = 8'd12;
        rom[374][51] = 8'd3;
        rom[374][52] = 8'd2;
        rom[374][53] = -8'd4;
        rom[374][54] = -8'd11;
        rom[374][55] = -8'd7;
        rom[374][56] = -8'd5;
        rom[374][57] = -8'd5;
        rom[374][58] = 8'd9;
        rom[374][59] = -8'd1;
        rom[374][60] = 8'd6;
        rom[374][61] = -8'd6;
        rom[374][62] = -8'd2;
        rom[374][63] = 8'd3;
        rom[375][0] = -8'd29;
        rom[375][1] = -8'd19;
        rom[375][2] = -8'd44;
        rom[375][3] = 8'd46;
        rom[375][4] = 8'd41;
        rom[375][5] = 8'd25;
        rom[375][6] = 8'd0;
        rom[375][7] = -8'd12;
        rom[375][8] = -8'd8;
        rom[375][9] = -8'd34;
        rom[375][10] = -8'd77;
        rom[375][11] = -8'd31;
        rom[375][12] = 8'd9;
        rom[375][13] = 8'd6;
        rom[375][14] = 8'd34;
        rom[375][15] = -8'd12;
        rom[375][16] = 8'd0;
        rom[375][17] = 8'd19;
        rom[375][18] = -8'd48;
        rom[375][19] = -8'd43;
        rom[375][20] = -8'd9;
        rom[375][21] = 8'd24;
        rom[375][22] = -8'd48;
        rom[375][23] = -8'd42;
        rom[375][24] = -8'd10;
        rom[375][25] = -8'd5;
        rom[375][26] = -8'd71;
        rom[375][27] = 8'd3;
        rom[375][28] = -8'd50;
        rom[375][29] = 8'd51;
        rom[375][30] = 8'd4;
        rom[375][31] = -8'd3;
        rom[375][32] = -8'd48;
        rom[375][33] = 8'd19;
        rom[375][34] = -8'd24;
        rom[375][35] = 8'd10;
        rom[375][36] = -8'd21;
        rom[375][37] = 8'd10;
        rom[375][38] = -8'd1;
        rom[375][39] = 8'd32;
        rom[375][40] = 8'd29;
        rom[375][41] = -8'd11;
        rom[375][42] = -8'd37;
        rom[375][43] = 8'd23;
        rom[375][44] = 8'd2;
        rom[375][45] = -8'd27;
        rom[375][46] = 8'd25;
        rom[375][47] = -8'd33;
        rom[375][48] = -8'd34;
        rom[375][49] = 8'd32;
        rom[375][50] = 8'd12;
        rom[375][51] = 8'd8;
        rom[375][52] = 8'd18;
        rom[375][53] = 8'd9;
        rom[375][54] = -8'd1;
        rom[375][55] = -8'd27;
        rom[375][56] = -8'd71;
        rom[375][57] = 8'd4;
        rom[375][58] = -8'd6;
        rom[375][59] = 8'd7;
        rom[375][60] = -8'd46;
        rom[375][61] = 8'd24;
        rom[375][62] = -8'd12;
        rom[375][63] = -8'd7;
        rom[376][0] = -8'd63;
        rom[376][1] = -8'd8;
        rom[376][2] = -8'd64;
        rom[376][3] = -8'd39;
        rom[376][4] = -8'd22;
        rom[376][5] = -8'd35;
        rom[376][6] = -8'd75;
        rom[376][7] = -8'd17;
        rom[376][8] = -8'd29;
        rom[376][9] = -8'd37;
        rom[376][10] = -8'd21;
        rom[376][11] = -8'd21;
        rom[376][12] = 8'd12;
        rom[376][13] = 8'd0;
        rom[376][14] = 8'd0;
        rom[376][15] = -8'd36;
        rom[376][16] = 8'd8;
        rom[376][17] = 8'd2;
        rom[376][18] = -8'd13;
        rom[376][19] = -8'd14;
        rom[376][20] = -8'd5;
        rom[376][21] = 8'd3;
        rom[376][22] = -8'd19;
        rom[376][23] = -8'd28;
        rom[376][24] = 8'd33;
        rom[376][25] = -8'd7;
        rom[376][26] = -8'd56;
        rom[376][27] = 8'd17;
        rom[376][28] = -8'd22;
        rom[376][29] = 8'd2;
        rom[376][30] = 8'd9;
        rom[376][31] = -8'd11;
        rom[376][32] = 8'd14;
        rom[376][33] = -8'd73;
        rom[376][34] = -8'd15;
        rom[376][35] = -8'd1;
        rom[376][36] = 8'd19;
        rom[376][37] = 8'd18;
        rom[376][38] = -8'd21;
        rom[376][39] = -8'd34;
        rom[376][40] = 8'd1;
        rom[376][41] = 8'd19;
        rom[376][42] = -8'd18;
        rom[376][43] = -8'd13;
        rom[376][44] = -8'd7;
        rom[376][45] = -8'd25;
        rom[376][46] = 8'd26;
        rom[376][47] = -8'd8;
        rom[376][48] = -8'd27;
        rom[376][49] = -8'd20;
        rom[376][50] = -8'd30;
        rom[376][51] = -8'd44;
        rom[376][52] = 8'd40;
        rom[376][53] = 8'd14;
        rom[376][54] = 8'd34;
        rom[376][55] = 8'd8;
        rom[376][56] = -8'd77;
        rom[376][57] = 8'd5;
        rom[376][58] = -8'd20;
        rom[376][59] = 8'd23;
        rom[376][60] = -8'd26;
        rom[376][61] = 8'd0;
        rom[376][62] = 8'd10;
        rom[376][63] = 8'd14;
        rom[377][0] = -8'd43;
        rom[377][1] = -8'd4;
        rom[377][2] = 8'd31;
        rom[377][3] = 8'd35;
        rom[377][4] = 8'd37;
        rom[377][5] = 8'd16;
        rom[377][6] = 8'd17;
        rom[377][7] = 8'd3;
        rom[377][8] = -8'd40;
        rom[377][9] = 8'd40;
        rom[377][10] = -8'd44;
        rom[377][11] = -8'd8;
        rom[377][12] = 8'd7;
        rom[377][13] = 8'd15;
        rom[377][14] = 8'd2;
        rom[377][15] = 8'd19;
        rom[377][16] = -8'd10;
        rom[377][17] = 8'd40;
        rom[377][18] = 8'd23;
        rom[377][19] = 8'd27;
        rom[377][20] = -8'd8;
        rom[377][21] = -8'd2;
        rom[377][22] = -8'd33;
        rom[377][23] = 8'd2;
        rom[377][24] = 8'd41;
        rom[377][25] = 8'd30;
        rom[377][26] = 8'd19;
        rom[377][27] = 8'd15;
        rom[377][28] = 8'd15;
        rom[377][29] = 8'd13;
        rom[377][30] = 8'd39;
        rom[377][31] = 8'd27;
        rom[377][32] = -8'd41;
        rom[377][33] = -8'd25;
        rom[377][34] = 8'd63;
        rom[377][35] = -8'd14;
        rom[377][36] = 8'd20;
        rom[377][37] = -8'd23;
        rom[377][38] = -8'd15;
        rom[377][39] = -8'd14;
        rom[377][40] = -8'd9;
        rom[377][41] = 8'd5;
        rom[377][42] = 8'd13;
        rom[377][43] = -8'd18;
        rom[377][44] = 8'd40;
        rom[377][45] = 8'd27;
        rom[377][46] = -8'd15;
        rom[377][47] = 8'd19;
        rom[377][48] = -8'd6;
        rom[377][49] = -8'd3;
        rom[377][50] = 8'd0;
        rom[377][51] = -8'd2;
        rom[377][52] = 8'd15;
        rom[377][53] = -8'd25;
        rom[377][54] = 8'd35;
        rom[377][55] = 8'd16;
        rom[377][56] = -8'd19;
        rom[377][57] = -8'd16;
        rom[377][58] = 8'd2;
        rom[377][59] = 8'd3;
        rom[377][60] = 8'd8;
        rom[377][61] = 8'd29;
        rom[377][62] = -8'd44;
        rom[377][63] = -8'd5;
        rom[378][0] = -8'd23;
        rom[378][1] = -8'd23;
        rom[378][2] = 8'd33;
        rom[378][3] = 8'd10;
        rom[378][4] = -8'd23;
        rom[378][5] = -8'd42;
        rom[378][6] = -8'd16;
        rom[378][7] = 8'd19;
        rom[378][8] = -8'd32;
        rom[378][9] = -8'd19;
        rom[378][10] = 8'd2;
        rom[378][11] = 8'd16;
        rom[378][12] = -8'd31;
        rom[378][13] = -8'd17;
        rom[378][14] = -8'd4;
        rom[378][15] = 8'd27;
        rom[378][16] = -8'd30;
        rom[378][17] = 8'd5;
        rom[378][18] = -8'd41;
        rom[378][19] = -8'd11;
        rom[378][20] = -8'd3;
        rom[378][21] = 8'd64;
        rom[378][22] = 8'd38;
        rom[378][23] = -8'd19;
        rom[378][24] = 8'd14;
        rom[378][25] = -8'd1;
        rom[378][26] = 8'd4;
        rom[378][27] = 8'd10;
        rom[378][28] = 8'd19;
        rom[378][29] = -8'd31;
        rom[378][30] = 8'd69;
        rom[378][31] = -8'd45;
        rom[378][32] = 8'd27;
        rom[378][33] = -8'd12;
        rom[378][34] = 8'd30;
        rom[378][35] = -8'd8;
        rom[378][36] = -8'd11;
        rom[378][37] = 8'd39;
        rom[378][38] = -8'd27;
        rom[378][39] = -8'd57;
        rom[378][40] = -8'd4;
        rom[378][41] = -8'd27;
        rom[378][42] = -8'd21;
        rom[378][43] = 8'd16;
        rom[378][44] = 8'd13;
        rom[378][45] = -8'd109;
        rom[378][46] = 8'd12;
        rom[378][47] = -8'd35;
        rom[378][48] = 8'd25;
        rom[378][49] = 8'd56;
        rom[378][50] = -8'd24;
        rom[378][51] = 8'd58;
        rom[378][52] = -8'd14;
        rom[378][53] = 8'd10;
        rom[378][54] = 8'd40;
        rom[378][55] = -8'd1;
        rom[378][56] = 8'd32;
        rom[378][57] = -8'd60;
        rom[378][58] = 8'd43;
        rom[378][59] = -8'd45;
        rom[378][60] = 8'd41;
        rom[378][61] = -8'd25;
        rom[378][62] = -8'd35;
        rom[378][63] = -8'd16;
        rom[379][0] = -8'd5;
        rom[379][1] = -8'd32;
        rom[379][2] = -8'd5;
        rom[379][3] = 8'd15;
        rom[379][4] = -8'd26;
        rom[379][5] = -8'd2;
        rom[379][6] = -8'd70;
        rom[379][7] = -8'd7;
        rom[379][8] = -8'd50;
        rom[379][9] = -8'd13;
        rom[379][10] = -8'd47;
        rom[379][11] = 8'd19;
        rom[379][12] = 8'd22;
        rom[379][13] = -8'd13;
        rom[379][14] = 8'd20;
        rom[379][15] = 8'd8;
        rom[379][16] = 8'd40;
        rom[379][17] = 8'd4;
        rom[379][18] = -8'd7;
        rom[379][19] = -8'd21;
        rom[379][20] = -8'd10;
        rom[379][21] = -8'd15;
        rom[379][22] = -8'd60;
        rom[379][23] = -8'd2;
        rom[379][24] = -8'd29;
        rom[379][25] = -8'd36;
        rom[379][26] = 8'd6;
        rom[379][27] = 8'd20;
        rom[379][28] = 8'd27;
        rom[379][29] = 8'd42;
        rom[379][30] = -8'd6;
        rom[379][31] = -8'd31;
        rom[379][32] = 8'd15;
        rom[379][33] = 8'd15;
        rom[379][34] = -8'd26;
        rom[379][35] = -8'd9;
        rom[379][36] = -8'd8;
        rom[379][37] = 8'd6;
        rom[379][38] = -8'd21;
        rom[379][39] = -8'd16;
        rom[379][40] = 8'd21;
        rom[379][41] = 8'd26;
        rom[379][42] = -8'd9;
        rom[379][43] = -8'd27;
        rom[379][44] = -8'd2;
        rom[379][45] = 8'd35;
        rom[379][46] = 8'd10;
        rom[379][47] = -8'd5;
        rom[379][48] = 8'd28;
        rom[379][49] = -8'd18;
        rom[379][50] = -8'd2;
        rom[379][51] = 8'd17;
        rom[379][52] = -8'd53;
        rom[379][53] = -8'd17;
        rom[379][54] = -8'd12;
        rom[379][55] = 8'd2;
        rom[379][56] = -8'd34;
        rom[379][57] = -8'd13;
        rom[379][58] = 8'd21;
        rom[379][59] = -8'd41;
        rom[379][60] = -8'd95;
        rom[379][61] = 8'd12;
        rom[379][62] = -8'd13;
        rom[379][63] = 8'd10;
        rom[380][0] = -8'd8;
        rom[380][1] = 8'd4;
        rom[380][2] = -8'd47;
        rom[380][3] = -8'd33;
        rom[380][4] = 8'd30;
        rom[380][5] = -8'd21;
        rom[380][6] = -8'd18;
        rom[380][7] = 8'd0;
        rom[380][8] = 8'd9;
        rom[380][9] = -8'd21;
        rom[380][10] = 8'd12;
        rom[380][11] = -8'd10;
        rom[380][12] = 8'd38;
        rom[380][13] = -8'd37;
        rom[380][14] = 8'd17;
        rom[380][15] = 8'd40;
        rom[380][16] = -8'd18;
        rom[380][17] = -8'd8;
        rom[380][18] = -8'd9;
        rom[380][19] = -8'd8;
        rom[380][20] = -8'd7;
        rom[380][21] = -8'd49;
        rom[380][22] = 8'd0;
        rom[380][23] = 8'd43;
        rom[380][24] = -8'd26;
        rom[380][25] = -8'd19;
        rom[380][26] = -8'd14;
        rom[380][27] = -8'd3;
        rom[380][28] = 8'd36;
        rom[380][29] = 8'd35;
        rom[380][30] = 8'd10;
        rom[380][31] = -8'd38;
        rom[380][32] = 8'd31;
        rom[380][33] = 8'd25;
        rom[380][34] = -8'd14;
        rom[380][35] = -8'd35;
        rom[380][36] = -8'd11;
        rom[380][37] = 8'd24;
        rom[380][38] = -8'd31;
        rom[380][39] = 8'd26;
        rom[380][40] = -8'd37;
        rom[380][41] = -8'd26;
        rom[380][42] = -8'd37;
        rom[380][43] = 8'd32;
        rom[380][44] = -8'd18;
        rom[380][45] = 8'd35;
        rom[380][46] = -8'd35;
        rom[380][47] = -8'd20;
        rom[380][48] = 8'd17;
        rom[380][49] = 8'd7;
        rom[380][50] = -8'd9;
        rom[380][51] = -8'd33;
        rom[380][52] = -8'd54;
        rom[380][53] = -8'd20;
        rom[380][54] = -8'd49;
        rom[380][55] = 8'd7;
        rom[380][56] = 8'd13;
        rom[380][57] = -8'd13;
        rom[380][58] = 8'd1;
        rom[380][59] = -8'd13;
        rom[380][60] = -8'd13;
        rom[380][61] = -8'd8;
        rom[380][62] = 8'd22;
        rom[380][63] = 8'd25;
        rom[381][0] = 8'd14;
        rom[381][1] = 8'd8;
        rom[381][2] = 8'd33;
        rom[381][3] = -8'd38;
        rom[381][4] = -8'd34;
        rom[381][5] = 8'd13;
        rom[381][6] = 8'd3;
        rom[381][7] = 8'd2;
        rom[381][8] = -8'd42;
        rom[381][9] = -8'd4;
        rom[381][10] = -8'd18;
        rom[381][11] = 8'd8;
        rom[381][12] = 8'd20;
        rom[381][13] = 8'd15;
        rom[381][14] = -8'd17;
        rom[381][15] = -8'd9;
        rom[381][16] = -8'd2;
        rom[381][17] = -8'd27;
        rom[381][18] = 8'd63;
        rom[381][19] = 8'd8;
        rom[381][20] = 8'd3;
        rom[381][21] = 8'd65;
        rom[381][22] = 8'd16;
        rom[381][23] = -8'd29;
        rom[381][24] = 8'd18;
        rom[381][25] = -8'd38;
        rom[381][26] = -8'd59;
        rom[381][27] = 8'd2;
        rom[381][28] = -8'd21;
        rom[381][29] = 8'd2;
        rom[381][30] = -8'd9;
        rom[381][31] = -8'd23;
        rom[381][32] = 8'd4;
        rom[381][33] = 8'd20;
        rom[381][34] = 8'd37;
        rom[381][35] = -8'd5;
        rom[381][36] = 8'd9;
        rom[381][37] = 8'd8;
        rom[381][38] = -8'd5;
        rom[381][39] = 8'd1;
        rom[381][40] = -8'd13;
        rom[381][41] = 8'd54;
        rom[381][42] = 8'd15;
        rom[381][43] = 8'd14;
        rom[381][44] = 8'd33;
        rom[381][45] = -8'd12;
        rom[381][46] = 8'd2;
        rom[381][47] = 8'd37;
        rom[381][48] = -8'd39;
        rom[381][49] = 8'd32;
        rom[381][50] = 8'd13;
        rom[381][51] = -8'd14;
        rom[381][52] = 8'd2;
        rom[381][53] = -8'd11;
        rom[381][54] = -8'd1;
        rom[381][55] = 8'd46;
        rom[381][56] = -8'd46;
        rom[381][57] = -8'd11;
        rom[381][58] = -8'd36;
        rom[381][59] = -8'd3;
        rom[381][60] = 8'd63;
        rom[381][61] = -8'd43;
        rom[381][62] = 8'd28;
        rom[381][63] = 8'd25;
        rom[382][0] = -8'd9;
        rom[382][1] = -8'd11;
        rom[382][2] = -8'd8;
        rom[382][3] = -8'd46;
        rom[382][4] = -8'd8;
        rom[382][5] = -8'd21;
        rom[382][6] = -8'd55;
        rom[382][7] = 8'd14;
        rom[382][8] = 8'd18;
        rom[382][9] = 8'd12;
        rom[382][10] = -8'd29;
        rom[382][11] = 8'd2;
        rom[382][12] = -8'd54;
        rom[382][13] = 8'd10;
        rom[382][14] = 8'd15;
        rom[382][15] = 8'd21;
        rom[382][16] = 8'd9;
        rom[382][17] = -8'd5;
        rom[382][18] = 8'd21;
        rom[382][19] = -8'd9;
        rom[382][20] = -8'd8;
        rom[382][21] = 8'd7;
        rom[382][22] = -8'd12;
        rom[382][23] = -8'd16;
        rom[382][24] = -8'd54;
        rom[382][25] = 8'd30;
        rom[382][26] = -8'd12;
        rom[382][27] = -8'd29;
        rom[382][28] = -8'd2;
        rom[382][29] = -8'd12;
        rom[382][30] = -8'd59;
        rom[382][31] = -8'd26;
        rom[382][32] = -8'd47;
        rom[382][33] = -8'd10;
        rom[382][34] = 8'd42;
        rom[382][35] = 8'd25;
        rom[382][36] = 8'd31;
        rom[382][37] = -8'd7;
        rom[382][38] = 8'd29;
        rom[382][39] = -8'd16;
        rom[382][40] = -8'd37;
        rom[382][41] = 8'd28;
        rom[382][42] = 8'd6;
        rom[382][43] = -8'd75;
        rom[382][44] = -8'd16;
        rom[382][45] = 8'd14;
        rom[382][46] = 8'd0;
        rom[382][47] = 8'd11;
        rom[382][48] = -8'd9;
        rom[382][49] = -8'd34;
        rom[382][50] = 8'd36;
        rom[382][51] = -8'd33;
        rom[382][52] = 8'd17;
        rom[382][53] = 8'd32;
        rom[382][54] = -8'd35;
        rom[382][55] = 8'd26;
        rom[382][56] = -8'd31;
        rom[382][57] = 8'd8;
        rom[382][58] = -8'd17;
        rom[382][59] = 8'd2;
        rom[382][60] = -8'd12;
        rom[382][61] = -8'd80;
        rom[382][62] = -8'd17;
        rom[382][63] = -8'd30;
        rom[383][0] = 8'd11;
        rom[383][1] = 8'd9;
        rom[383][2] = 8'd31;
        rom[383][3] = -8'd36;
        rom[383][4] = -8'd17;
        rom[383][5] = -8'd16;
        rom[383][6] = 8'd18;
        rom[383][7] = -8'd6;
        rom[383][8] = -8'd39;
        rom[383][9] = -8'd53;
        rom[383][10] = -8'd15;
        rom[383][11] = 8'd5;
        rom[383][12] = -8'd34;
        rom[383][13] = 8'd5;
        rom[383][14] = 8'd35;
        rom[383][15] = 8'd3;
        rom[383][16] = -8'd20;
        rom[383][17] = 8'd17;
        rom[383][18] = 8'd3;
        rom[383][19] = -8'd9;
        rom[383][20] = -8'd6;
        rom[383][21] = -8'd6;
        rom[383][22] = 8'd23;
        rom[383][23] = 8'd29;
        rom[383][24] = -8'd49;
        rom[383][25] = 8'd48;
        rom[383][26] = -8'd21;
        rom[383][27] = 8'd25;
        rom[383][28] = -8'd22;
        rom[383][29] = 8'd8;
        rom[383][30] = 8'd12;
        rom[383][31] = -8'd22;
        rom[383][32] = 8'd17;
        rom[383][33] = 8'd32;
        rom[383][34] = -8'd14;
        rom[383][35] = -8'd24;
        rom[383][36] = 8'd3;
        rom[383][37] = 8'd0;
        rom[383][38] = 8'd35;
        rom[383][39] = 8'd8;
        rom[383][40] = 8'd25;
        rom[383][41] = 8'd3;
        rom[383][42] = -8'd18;
        rom[383][43] = 8'd7;
        rom[383][44] = 8'd2;
        rom[383][45] = -8'd30;
        rom[383][46] = 8'd1;
        rom[383][47] = -8'd37;
        rom[383][48] = 8'd15;
        rom[383][49] = -8'd9;
        rom[383][50] = -8'd9;
        rom[383][51] = -8'd49;
        rom[383][52] = 8'd24;
        rom[383][53] = 8'd13;
        rom[383][54] = 8'd5;
        rom[383][55] = -8'd18;
        rom[383][56] = 8'd52;
        rom[383][57] = -8'd34;
        rom[383][58] = 8'd13;
        rom[383][59] = -8'd51;
        rom[383][60] = 8'd15;
        rom[383][61] = -8'd32;
        rom[383][62] = -8'd49;
        rom[383][63] = 8'd6;
        rom[384][0] = -8'd3;
        rom[384][1] = 8'd6;
        rom[384][2] = -8'd5;
        rom[384][3] = -8'd3;
        rom[384][4] = -8'd42;
        rom[384][5] = 8'd26;
        rom[384][6] = -8'd3;
        rom[384][7] = 8'd7;
        rom[384][8] = -8'd40;
        rom[384][9] = 8'd3;
        rom[384][10] = 8'd29;
        rom[384][11] = 8'd1;
        rom[384][12] = 8'd0;
        rom[384][13] = -8'd14;
        rom[384][14] = -8'd33;
        rom[384][15] = -8'd15;
        rom[384][16] = 8'd15;
        rom[384][17] = 8'd24;
        rom[384][18] = 8'd5;
        rom[384][19] = -8'd16;
        rom[384][20] = -8'd3;
        rom[384][21] = -8'd4;
        rom[384][22] = -8'd18;
        rom[384][23] = 8'd6;
        rom[384][24] = -8'd20;
        rom[384][25] = -8'd18;
        rom[384][26] = 8'd20;
        rom[384][27] = -8'd23;
        rom[384][28] = 8'd7;
        rom[384][29] = 8'd11;
        rom[384][30] = -8'd22;
        rom[384][31] = 8'd8;
        rom[384][32] = -8'd40;
        rom[384][33] = 8'd14;
        rom[384][34] = -8'd1;
        rom[384][35] = -8'd40;
        rom[384][36] = -8'd7;
        rom[384][37] = -8'd23;
        rom[384][38] = -8'd4;
        rom[384][39] = 8'd24;
        rom[384][40] = -8'd52;
        rom[384][41] = -8'd38;
        rom[384][42] = -8'd4;
        rom[384][43] = -8'd18;
        rom[384][44] = -8'd62;
        rom[384][45] = 8'd7;
        rom[384][46] = 8'd6;
        rom[384][47] = -8'd38;
        rom[384][48] = -8'd49;
        rom[384][49] = -8'd39;
        rom[384][50] = -8'd1;
        rom[384][51] = -8'd43;
        rom[384][52] = 8'd30;
        rom[384][53] = -8'd27;
        rom[384][54] = 8'd9;
        rom[384][55] = 8'd1;
        rom[384][56] = 8'd5;
        rom[384][57] = 8'd18;
        rom[384][58] = -8'd22;
        rom[384][59] = 8'd9;
        rom[384][60] = 8'd3;
        rom[384][61] = -8'd30;
        rom[384][62] = -8'd38;
        rom[384][63] = 8'd26;
        rom[385][0] = -8'd5;
        rom[385][1] = -8'd35;
        rom[385][2] = 8'd41;
        rom[385][3] = -8'd34;
        rom[385][4] = -8'd48;
        rom[385][5] = 8'd60;
        rom[385][6] = -8'd94;
        rom[385][7] = -8'd20;
        rom[385][8] = 8'd24;
        rom[385][9] = -8'd32;
        rom[385][10] = -8'd17;
        rom[385][11] = -8'd24;
        rom[385][12] = 8'd49;
        rom[385][13] = -8'd7;
        rom[385][14] = 8'd23;
        rom[385][15] = 8'd20;
        rom[385][16] = -8'd28;
        rom[385][17] = 8'd2;
        rom[385][18] = -8'd21;
        rom[385][19] = 8'd31;
        rom[385][20] = -8'd6;
        rom[385][21] = 8'd23;
        rom[385][22] = -8'd7;
        rom[385][23] = -8'd11;
        rom[385][24] = 8'd1;
        rom[385][25] = 8'd11;
        rom[385][26] = -8'd8;
        rom[385][27] = -8'd14;
        rom[385][28] = 8'd14;
        rom[385][29] = -8'd42;
        rom[385][30] = 8'd16;
        rom[385][31] = -8'd4;
        rom[385][32] = 8'd37;
        rom[385][33] = 8'd4;
        rom[385][34] = 8'd19;
        rom[385][35] = -8'd22;
        rom[385][36] = -8'd3;
        rom[385][37] = -8'd15;
        rom[385][38] = 8'd25;
        rom[385][39] = 8'd29;
        rom[385][40] = 8'd47;
        rom[385][41] = -8'd12;
        rom[385][42] = 8'd29;
        rom[385][43] = -8'd13;
        rom[385][44] = -8'd16;
        rom[385][45] = 8'd21;
        rom[385][46] = -8'd7;
        rom[385][47] = 8'd43;
        rom[385][48] = -8'd3;
        rom[385][49] = 8'd43;
        rom[385][50] = 8'd4;
        rom[385][51] = 8'd4;
        rom[385][52] = -8'd52;
        rom[385][53] = -8'd13;
        rom[385][54] = -8'd15;
        rom[385][55] = 8'd10;
        rom[385][56] = 8'd34;
        rom[385][57] = 8'd10;
        rom[385][58] = -8'd66;
        rom[385][59] = -8'd2;
        rom[385][60] = -8'd58;
        rom[385][61] = 8'd13;
        rom[385][62] = -8'd33;
        rom[385][63] = -8'd10;
        rom[386][0] = 8'd30;
        rom[386][1] = 8'd25;
        rom[386][2] = -8'd51;
        rom[386][3] = -8'd16;
        rom[386][4] = -8'd69;
        rom[386][5] = 8'd1;
        rom[386][6] = -8'd119;
        rom[386][7] = 8'd2;
        rom[386][8] = -8'd57;
        rom[386][9] = -8'd16;
        rom[386][10] = 8'd53;
        rom[386][11] = -8'd5;
        rom[386][12] = -8'd5;
        rom[386][13] = -8'd58;
        rom[386][14] = -8'd77;
        rom[386][15] = 8'd20;
        rom[386][16] = 8'd43;
        rom[386][17] = -8'd15;
        rom[386][18] = 8'd12;
        rom[386][19] = -8'd32;
        rom[386][20] = -8'd10;
        rom[386][21] = 8'd53;
        rom[386][22] = -8'd41;
        rom[386][23] = 8'd11;
        rom[386][24] = -8'd74;
        rom[386][25] = -8'd2;
        rom[386][26] = 8'd21;
        rom[386][27] = -8'd11;
        rom[386][28] = -8'd3;
        rom[386][29] = -8'd16;
        rom[386][30] = 8'd28;
        rom[386][31] = -8'd34;
        rom[386][32] = 8'd29;
        rom[386][33] = -8'd78;
        rom[386][34] = -8'd11;
        rom[386][35] = -8'd40;
        rom[386][36] = -8'd63;
        rom[386][37] = -8'd4;
        rom[386][38] = 8'd11;
        rom[386][39] = -8'd20;
        rom[386][40] = -8'd4;
        rom[386][41] = 8'd24;
        rom[386][42] = -8'd65;
        rom[386][43] = -8'd20;
        rom[386][44] = 8'd4;
        rom[386][45] = -8'd31;
        rom[386][46] = 8'd67;
        rom[386][47] = 8'd6;
        rom[386][48] = 8'd15;
        rom[386][49] = -8'd25;
        rom[386][50] = 8'd3;
        rom[386][51] = -8'd32;
        rom[386][52] = -8'd35;
        rom[386][53] = -8'd55;
        rom[386][54] = -8'd8;
        rom[386][55] = -8'd3;
        rom[386][56] = -8'd20;
        rom[386][57] = 8'd5;
        rom[386][58] = -8'd21;
        rom[386][59] = -8'd8;
        rom[386][60] = -8'd9;
        rom[386][61] = 8'd18;
        rom[386][62] = -8'd21;
        rom[386][63] = 8'd6;
        rom[387][0] = -8'd12;
        rom[387][1] = 8'd8;
        rom[387][2] = -8'd12;
        rom[387][3] = 8'd18;
        rom[387][4] = 8'd13;
        rom[387][5] = 8'd15;
        rom[387][6] = 8'd5;
        rom[387][7] = 8'd33;
        rom[387][8] = 8'd9;
        rom[387][9] = 8'd15;
        rom[387][10] = 8'd25;
        rom[387][11] = -8'd17;
        rom[387][12] = -8'd26;
        rom[387][13] = -8'd44;
        rom[387][14] = 8'd28;
        rom[387][15] = 8'd26;
        rom[387][16] = -8'd24;
        rom[387][17] = 8'd11;
        rom[387][18] = 8'd17;
        rom[387][19] = -8'd38;
        rom[387][20] = 8'd1;
        rom[387][21] = -8'd7;
        rom[387][22] = 8'd5;
        rom[387][23] = -8'd6;
        rom[387][24] = -8'd29;
        rom[387][25] = -8'd46;
        rom[387][26] = 8'd39;
        rom[387][27] = 8'd12;
        rom[387][28] = 8'd8;
        rom[387][29] = 8'd30;
        rom[387][30] = 8'd8;
        rom[387][31] = 8'd16;
        rom[387][32] = -8'd42;
        rom[387][33] = -8'd33;
        rom[387][34] = 8'd15;
        rom[387][35] = 8'd1;
        rom[387][36] = 8'd5;
        rom[387][37] = 8'd43;
        rom[387][38] = -8'd60;
        rom[387][39] = 8'd23;
        rom[387][40] = -8'd10;
        rom[387][41] = 8'd38;
        rom[387][42] = 8'd19;
        rom[387][43] = -8'd8;
        rom[387][44] = 8'd30;
        rom[387][45] = -8'd31;
        rom[387][46] = -8'd41;
        rom[387][47] = -8'd30;
        rom[387][48] = 8'd0;
        rom[387][49] = -8'd31;
        rom[387][50] = -8'd4;
        rom[387][51] = 8'd3;
        rom[387][52] = 8'd54;
        rom[387][53] = -8'd44;
        rom[387][54] = -8'd22;
        rom[387][55] = -8'd31;
        rom[387][56] = -8'd7;
        rom[387][57] = -8'd42;
        rom[387][58] = 8'd33;
        rom[387][59] = -8'd25;
        rom[387][60] = 8'd23;
        rom[387][61] = -8'd63;
        rom[387][62] = 8'd18;
        rom[387][63] = 8'd16;
        rom[388][0] = 8'd19;
        rom[388][1] = -8'd53;
        rom[388][2] = -8'd14;
        rom[388][3] = -8'd21;
        rom[388][4] = 8'd11;
        rom[388][5] = -8'd17;
        rom[388][6] = -8'd10;
        rom[388][7] = 8'd27;
        rom[388][8] = -8'd18;
        rom[388][9] = -8'd18;
        rom[388][10] = -8'd39;
        rom[388][11] = 8'd22;
        rom[388][12] = 8'd3;
        rom[388][13] = -8'd17;
        rom[388][14] = -8'd26;
        rom[388][15] = -8'd22;
        rom[388][16] = -8'd2;
        rom[388][17] = -8'd16;
        rom[388][18] = -8'd32;
        rom[388][19] = 8'd32;
        rom[388][20] = -8'd14;
        rom[388][21] = 8'd7;
        rom[388][22] = -8'd38;
        rom[388][23] = -8'd9;
        rom[388][24] = 8'd14;
        rom[388][25] = -8'd37;
        rom[388][26] = -8'd25;
        rom[388][27] = 8'd12;
        rom[388][28] = 8'd3;
        rom[388][29] = -8'd28;
        rom[388][30] = -8'd5;
        rom[388][31] = -8'd24;
        rom[388][32] = 8'd38;
        rom[388][33] = -8'd12;
        rom[388][34] = 8'd4;
        rom[388][35] = 8'd3;
        rom[388][36] = -8'd24;
        rom[388][37] = -8'd11;
        rom[388][38] = -8'd26;
        rom[388][39] = -8'd42;
        rom[388][40] = 8'd28;
        rom[388][41] = -8'd13;
        rom[388][42] = -8'd21;
        rom[388][43] = -8'd19;
        rom[388][44] = -8'd7;
        rom[388][45] = 8'd22;
        rom[388][46] = -8'd11;
        rom[388][47] = -8'd54;
        rom[388][48] = 8'd28;
        rom[388][49] = -8'd16;
        rom[388][50] = -8'd3;
        rom[388][51] = -8'd7;
        rom[388][52] = -8'd2;
        rom[388][53] = -8'd40;
        rom[388][54] = 8'd2;
        rom[388][55] = -8'd56;
        rom[388][56] = -8'd13;
        rom[388][57] = 8'd37;
        rom[388][58] = 8'd15;
        rom[388][59] = -8'd43;
        rom[388][60] = 8'd28;
        rom[388][61] = -8'd5;
        rom[388][62] = 8'd6;
        rom[388][63] = -8'd42;
        rom[389][0] = -8'd1;
        rom[389][1] = 8'd2;
        rom[389][2] = 8'd3;
        rom[389][3] = 8'd5;
        rom[389][4] = -8'd4;
        rom[389][5] = -8'd6;
        rom[389][6] = -8'd3;
        rom[389][7] = -8'd1;
        rom[389][8] = 8'd7;
        rom[389][9] = -8'd5;
        rom[389][10] = 8'd10;
        rom[389][11] = 8'd2;
        rom[389][12] = -8'd9;
        rom[389][13] = -8'd2;
        rom[389][14] = 8'd5;
        rom[389][15] = -8'd1;
        rom[389][16] = 8'd12;
        rom[389][17] = 8'd7;
        rom[389][18] = -8'd4;
        rom[389][19] = -8'd3;
        rom[389][20] = -8'd6;
        rom[389][21] = -8'd1;
        rom[389][22] = 8'd5;
        rom[389][23] = 8'd7;
        rom[389][24] = 8'd22;
        rom[389][25] = 8'd3;
        rom[389][26] = 8'd4;
        rom[389][27] = -8'd9;
        rom[389][28] = -8'd12;
        rom[389][29] = -8'd5;
        rom[389][30] = 8'd1;
        rom[389][31] = 8'd5;
        rom[389][32] = -8'd8;
        rom[389][33] = 8'd5;
        rom[389][34] = 8'd0;
        rom[389][35] = 8'd11;
        rom[389][36] = 8'd11;
        rom[389][37] = -8'd2;
        rom[389][38] = -8'd4;
        rom[389][39] = -8'd4;
        rom[389][40] = -8'd9;
        rom[389][41] = 8'd6;
        rom[389][42] = 8'd6;
        rom[389][43] = 8'd2;
        rom[389][44] = -8'd6;
        rom[389][45] = 8'd4;
        rom[389][46] = -8'd1;
        rom[389][47] = -8'd13;
        rom[389][48] = 8'd1;
        rom[389][49] = -8'd10;
        rom[389][50] = 8'd3;
        rom[389][51] = 8'd1;
        rom[389][52] = 8'd4;
        rom[389][53] = 8'd3;
        rom[389][54] = 8'd2;
        rom[389][55] = 8'd7;
        rom[389][56] = 8'd0;
        rom[389][57] = 8'd0;
        rom[389][58] = 8'd2;
        rom[389][59] = -8'd4;
        rom[389][60] = -8'd8;
        rom[389][61] = 8'd8;
        rom[389][62] = 8'd8;
        rom[389][63] = -8'd3;
        rom[390][0] = 8'd9;
        rom[390][1] = -8'd11;
        rom[390][2] = -8'd3;
        rom[390][3] = -8'd11;
        rom[390][4] = -8'd57;
        rom[390][5] = 8'd24;
        rom[390][6] = -8'd40;
        rom[390][7] = -8'd25;
        rom[390][8] = 8'd15;
        rom[390][9] = 8'd17;
        rom[390][10] = -8'd24;
        rom[390][11] = 8'd34;
        rom[390][12] = 8'd7;
        rom[390][13] = 8'd9;
        rom[390][14] = -8'd82;
        rom[390][15] = -8'd16;
        rom[390][16] = -8'd10;
        rom[390][17] = 8'd34;
        rom[390][18] = 8'd21;
        rom[390][19] = -8'd37;
        rom[390][20] = -8'd3;
        rom[390][21] = -8'd24;
        rom[390][22] = 8'd9;
        rom[390][23] = 8'd32;
        rom[390][24] = -8'd11;
        rom[390][25] = -8'd1;
        rom[390][26] = 8'd17;
        rom[390][27] = 8'd16;
        rom[390][28] = -8'd14;
        rom[390][29] = 8'd29;
        rom[390][30] = -8'd17;
        rom[390][31] = 8'd41;
        rom[390][32] = 8'd0;
        rom[390][33] = -8'd20;
        rom[390][34] = 8'd18;
        rom[390][35] = 8'd4;
        rom[390][36] = -8'd24;
        rom[390][37] = 8'd10;
        rom[390][38] = 8'd19;
        rom[390][39] = -8'd26;
        rom[390][40] = 8'd27;
        rom[390][41] = 8'd3;
        rom[390][42] = 8'd3;
        rom[390][43] = 8'd3;
        rom[390][44] = 8'd44;
        rom[390][45] = 8'd15;
        rom[390][46] = 8'd10;
        rom[390][47] = -8'd21;
        rom[390][48] = -8'd15;
        rom[390][49] = -8'd37;
        rom[390][50] = 8'd15;
        rom[390][51] = 8'd8;
        rom[390][52] = -8'd34;
        rom[390][53] = -8'd48;
        rom[390][54] = 8'd10;
        rom[390][55] = 8'd29;
        rom[390][56] = 8'd46;
        rom[390][57] = 8'd19;
        rom[390][58] = 8'd24;
        rom[390][59] = -8'd8;
        rom[390][60] = -8'd10;
        rom[390][61] = -8'd50;
        rom[390][62] = -8'd6;
        rom[390][63] = 8'd21;
        rom[391][0] = 8'd63;
        rom[391][1] = 8'd41;
        rom[391][2] = 8'd8;
        rom[391][3] = -8'd35;
        rom[391][4] = 8'd0;
        rom[391][5] = -8'd15;
        rom[391][6] = 8'd19;
        rom[391][7] = 8'd55;
        rom[391][8] = 8'd19;
        rom[391][9] = -8'd10;
        rom[391][10] = 8'd10;
        rom[391][11] = -8'd46;
        rom[391][12] = -8'd94;
        rom[391][13] = 8'd43;
        rom[391][14] = -8'd11;
        rom[391][15] = 8'd39;
        rom[391][16] = -8'd31;
        rom[391][17] = -8'd35;
        rom[391][18] = 8'd24;
        rom[391][19] = 8'd63;
        rom[391][20] = -8'd5;
        rom[391][21] = 8'd14;
        rom[391][22] = 8'd19;
        rom[391][23] = 8'd10;
        rom[391][24] = 8'd34;
        rom[391][25] = -8'd29;
        rom[391][26] = -8'd13;
        rom[391][27] = -8'd28;
        rom[391][28] = 8'd7;
        rom[391][29] = -8'd43;
        rom[391][30] = -8'd15;
        rom[391][31] = -8'd123;
        rom[391][32] = 8'd45;
        rom[391][33] = 8'd28;
        rom[391][34] = 8'd50;
        rom[391][35] = 8'd42;
        rom[391][36] = -8'd5;
        rom[391][37] = 8'd51;
        rom[391][38] = 8'd1;
        rom[391][39] = -8'd10;
        rom[391][40] = -8'd19;
        rom[391][41] = -8'd7;
        rom[391][42] = 8'd22;
        rom[391][43] = 8'd7;
        rom[391][44] = 8'd17;
        rom[391][45] = 8'd44;
        rom[391][46] = -8'd11;
        rom[391][47] = -8'd2;
        rom[391][48] = 8'd31;
        rom[391][49] = 8'd2;
        rom[391][50] = 8'd6;
        rom[391][51] = -8'd18;
        rom[391][52] = 8'd7;
        rom[391][53] = 8'd21;
        rom[391][54] = 8'd30;
        rom[391][55] = -8'd14;
        rom[391][56] = 8'd24;
        rom[391][57] = -8'd7;
        rom[391][58] = -8'd26;
        rom[391][59] = -8'd16;
        rom[391][60] = -8'd13;
        rom[391][61] = -8'd8;
        rom[391][62] = -8'd13;
        rom[391][63] = 8'd33;
        rom[392][0] = 8'd19;
        rom[392][1] = 8'd8;
        rom[392][2] = -8'd26;
        rom[392][3] = -8'd11;
        rom[392][4] = 8'd21;
        rom[392][5] = -8'd44;
        rom[392][6] = -8'd14;
        rom[392][7] = -8'd60;
        rom[392][8] = -8'd2;
        rom[392][9] = -8'd26;
        rom[392][10] = -8'd23;
        rom[392][11] = -8'd3;
        rom[392][12] = -8'd13;
        rom[392][13] = -8'd24;
        rom[392][14] = 8'd38;
        rom[392][15] = 8'd0;
        rom[392][16] = -8'd19;
        rom[392][17] = -8'd29;
        rom[392][18] = 8'd31;
        rom[392][19] = -8'd1;
        rom[392][20] = 8'd5;
        rom[392][21] = -8'd23;
        rom[392][22] = 8'd17;
        rom[392][23] = -8'd18;
        rom[392][24] = -8'd10;
        rom[392][25] = 8'd4;
        rom[392][26] = -8'd35;
        rom[392][27] = -8'd30;
        rom[392][28] = -8'd3;
        rom[392][29] = 8'd19;
        rom[392][30] = -8'd75;
        rom[392][31] = 8'd3;
        rom[392][32] = -8'd6;
        rom[392][33] = 8'd6;
        rom[392][34] = -8'd14;
        rom[392][35] = 8'd12;
        rom[392][36] = -8'd3;
        rom[392][37] = -8'd41;
        rom[392][38] = -8'd42;
        rom[392][39] = 8'd7;
        rom[392][40] = -8'd36;
        rom[392][41] = -8'd5;
        rom[392][42] = -8'd93;
        rom[392][43] = 8'd17;
        rom[392][44] = -8'd36;
        rom[392][45] = -8'd20;
        rom[392][46] = -8'd14;
        rom[392][47] = -8'd23;
        rom[392][48] = -8'd10;
        rom[392][49] = 8'd12;
        rom[392][50] = 8'd3;
        rom[392][51] = -8'd35;
        rom[392][52] = 8'd60;
        rom[392][53] = -8'd1;
        rom[392][54] = -8'd46;
        rom[392][55] = 8'd45;
        rom[392][56] = 8'd10;
        rom[392][57] = 8'd14;
        rom[392][58] = -8'd3;
        rom[392][59] = -8'd12;
        rom[392][60] = -8'd1;
        rom[392][61] = 8'd6;
        rom[392][62] = -8'd21;
        rom[392][63] = 8'd9;
        rom[393][0] = -8'd27;
        rom[393][1] = -8'd51;
        rom[393][2] = 8'd2;
        rom[393][3] = -8'd55;
        rom[393][4] = -8'd13;
        rom[393][5] = 8'd19;
        rom[393][6] = -8'd3;
        rom[393][7] = 8'd11;
        rom[393][8] = -8'd46;
        rom[393][9] = 8'd14;
        rom[393][10] = 8'd3;
        rom[393][11] = 8'd22;
        rom[393][12] = -8'd3;
        rom[393][13] = -8'd22;
        rom[393][14] = -8'd2;
        rom[393][15] = -8'd45;
        rom[393][16] = 8'd0;
        rom[393][17] = -8'd23;
        rom[393][18] = -8'd19;
        rom[393][19] = -8'd46;
        rom[393][20] = -8'd1;
        rom[393][21] = -8'd8;
        rom[393][22] = 8'd2;
        rom[393][23] = -8'd13;
        rom[393][24] = 8'd22;
        rom[393][25] = 8'd3;
        rom[393][26] = 8'd9;
        rom[393][27] = -8'd1;
        rom[393][28] = 8'd36;
        rom[393][29] = -8'd7;
        rom[393][30] = -8'd25;
        rom[393][31] = 8'd21;
        rom[393][32] = -8'd3;
        rom[393][33] = -8'd32;
        rom[393][34] = 8'd11;
        rom[393][35] = -8'd27;
        rom[393][36] = -8'd10;
        rom[393][37] = -8'd16;
        rom[393][38] = -8'd27;
        rom[393][39] = 8'd9;
        rom[393][40] = 8'd19;
        rom[393][41] = -8'd6;
        rom[393][42] = -8'd44;
        rom[393][43] = -8'd4;
        rom[393][44] = -8'd11;
        rom[393][45] = -8'd12;
        rom[393][46] = -8'd28;
        rom[393][47] = 8'd17;
        rom[393][48] = -8'd10;
        rom[393][49] = -8'd28;
        rom[393][50] = -8'd57;
        rom[393][51] = 8'd13;
        rom[393][52] = -8'd2;
        rom[393][53] = 8'd16;
        rom[393][54] = -8'd29;
        rom[393][55] = 8'd21;
        rom[393][56] = 8'd3;
        rom[393][57] = 8'd33;
        rom[393][58] = 8'd31;
        rom[393][59] = -8'd21;
        rom[393][60] = -8'd35;
        rom[393][61] = -8'd4;
        rom[393][62] = 8'd37;
        rom[393][63] = 8'd57;
        rom[394][0] = -8'd5;
        rom[394][1] = -8'd51;
        rom[394][2] = 8'd11;
        rom[394][3] = 8'd40;
        rom[394][4] = -8'd21;
        rom[394][5] = -8'd33;
        rom[394][6] = -8'd7;
        rom[394][7] = -8'd30;
        rom[394][8] = -8'd8;
        rom[394][9] = -8'd21;
        rom[394][10] = -8'd2;
        rom[394][11] = -8'd15;
        rom[394][12] = 8'd10;
        rom[394][13] = 8'd10;
        rom[394][14] = -8'd52;
        rom[394][15] = 8'd46;
        rom[394][16] = -8'd21;
        rom[394][17] = -8'd61;
        rom[394][18] = -8'd68;
        rom[394][19] = -8'd4;
        rom[394][20] = -8'd13;
        rom[394][21] = -8'd39;
        rom[394][22] = 8'd44;
        rom[394][23] = -8'd24;
        rom[394][24] = -8'd18;
        rom[394][25] = -8'd3;
        rom[394][26] = -8'd7;
        rom[394][27] = -8'd10;
        rom[394][28] = -8'd33;
        rom[394][29] = -8'd35;
        rom[394][30] = 8'd33;
        rom[394][31] = -8'd49;
        rom[394][32] = 8'd24;
        rom[394][33] = -8'd18;
        rom[394][34] = -8'd36;
        rom[394][35] = 8'd29;
        rom[394][36] = -8'd49;
        rom[394][37] = 8'd71;
        rom[394][38] = -8'd4;
        rom[394][39] = -8'd44;
        rom[394][40] = -8'd16;
        rom[394][41] = -8'd33;
        rom[394][42] = 8'd31;
        rom[394][43] = -8'd5;
        rom[394][44] = 8'd21;
        rom[394][45] = -8'd16;
        rom[394][46] = 8'd11;
        rom[394][47] = 8'd38;
        rom[394][48] = 8'd20;
        rom[394][49] = 8'd12;
        rom[394][50] = -8'd26;
        rom[394][51] = 8'd2;
        rom[394][52] = -8'd15;
        rom[394][53] = -8'd50;
        rom[394][54] = -8'd15;
        rom[394][55] = -8'd4;
        rom[394][56] = 8'd27;
        rom[394][57] = -8'd7;
        rom[394][58] = 8'd6;
        rom[394][59] = 8'd27;
        rom[394][60] = 8'd41;
        rom[394][61] = 8'd1;
        rom[394][62] = 8'd30;
        rom[394][63] = -8'd29;
        rom[395][0] = -8'd39;
        rom[395][1] = 8'd14;
        rom[395][2] = 8'd0;
        rom[395][3] = -8'd37;
        rom[395][4] = 8'd23;
        rom[395][5] = -8'd4;
        rom[395][6] = 8'd9;
        rom[395][7] = -8'd57;
        rom[395][8] = -8'd2;
        rom[395][9] = -8'd9;
        rom[395][10] = -8'd52;
        rom[395][11] = -8'd4;
        rom[395][12] = 8'd3;
        rom[395][13] = 8'd21;
        rom[395][14] = -8'd12;
        rom[395][15] = -8'd11;
        rom[395][16] = -8'd22;
        rom[395][17] = -8'd12;
        rom[395][18] = -8'd46;
        rom[395][19] = -8'd8;
        rom[395][20] = -8'd8;
        rom[395][21] = 8'd12;
        rom[395][22] = -8'd9;
        rom[395][23] = -8'd3;
        rom[395][24] = -8'd7;
        rom[395][25] = -8'd3;
        rom[395][26] = -8'd4;
        rom[395][27] = -8'd20;
        rom[395][28] = -8'd36;
        rom[395][29] = -8'd82;
        rom[395][30] = -8'd19;
        rom[395][31] = -8'd18;
        rom[395][32] = 8'd3;
        rom[395][33] = 8'd11;
        rom[395][34] = 8'd46;
        rom[395][35] = 8'd47;
        rom[395][36] = -8'd14;
        rom[395][37] = -8'd69;
        rom[395][38] = -8'd47;
        rom[395][39] = -8'd42;
        rom[395][40] = -8'd1;
        rom[395][41] = 8'd12;
        rom[395][42] = 8'd21;
        rom[395][43] = 8'd20;
        rom[395][44] = -8'd8;
        rom[395][45] = 8'd0;
        rom[395][46] = 8'd26;
        rom[395][47] = -8'd15;
        rom[395][48] = -8'd59;
        rom[395][49] = 8'd28;
        rom[395][50] = -8'd10;
        rom[395][51] = 8'd9;
        rom[395][52] = 8'd5;
        rom[395][53] = -8'd29;
        rom[395][54] = -8'd1;
        rom[395][55] = -8'd53;
        rom[395][56] = 8'd1;
        rom[395][57] = 8'd2;
        rom[395][58] = -8'd26;
        rom[395][59] = -8'd9;
        rom[395][60] = 8'd6;
        rom[395][61] = 8'd7;
        rom[395][62] = -8'd14;
        rom[395][63] = -8'd19;
        rom[396][0] = -8'd73;
        rom[396][1] = -8'd49;
        rom[396][2] = -8'd54;
        rom[396][3] = 8'd13;
        rom[396][4] = 8'd34;
        rom[396][5] = 8'd14;
        rom[396][6] = -8'd38;
        rom[396][7] = -8'd5;
        rom[396][8] = -8'd8;
        rom[396][9] = -8'd26;
        rom[396][10] = 8'd1;
        rom[396][11] = 8'd39;
        rom[396][12] = -8'd49;
        rom[396][13] = -8'd58;
        rom[396][14] = 8'd8;
        rom[396][15] = 8'd4;
        rom[396][16] = -8'd16;
        rom[396][17] = -8'd15;
        rom[396][18] = 8'd31;
        rom[396][19] = -8'd15;
        rom[396][20] = -8'd3;
        rom[396][21] = -8'd19;
        rom[396][22] = 8'd50;
        rom[396][23] = -8'd5;
        rom[396][24] = 8'd18;
        rom[396][25] = -8'd2;
        rom[396][26] = 8'd18;
        rom[396][27] = -8'd14;
        rom[396][28] = 8'd31;
        rom[396][29] = 8'd16;
        rom[396][30] = 8'd51;
        rom[396][31] = -8'd20;
        rom[396][32] = 8'd23;
        rom[396][33] = 8'd37;
        rom[396][34] = 8'd23;
        rom[396][35] = 8'd35;
        rom[396][36] = -8'd8;
        rom[396][37] = 8'd11;
        rom[396][38] = 8'd1;
        rom[396][39] = 8'd44;
        rom[396][40] = -8'd55;
        rom[396][41] = 8'd19;
        rom[396][42] = 8'd5;
        rom[396][43] = 8'd56;
        rom[396][44] = -8'd9;
        rom[396][45] = 8'd36;
        rom[396][46] = 8'd20;
        rom[396][47] = -8'd17;
        rom[396][48] = -8'd4;
        rom[396][49] = 8'd8;
        rom[396][50] = 8'd25;
        rom[396][51] = 8'd3;
        rom[396][52] = 8'd18;
        rom[396][53] = -8'd7;
        rom[396][54] = 8'd45;
        rom[396][55] = 8'd1;
        rom[396][56] = -8'd24;
        rom[396][57] = -8'd47;
        rom[396][58] = -8'd27;
        rom[396][59] = -8'd20;
        rom[396][60] = 8'd10;
        rom[396][61] = 8'd9;
        rom[396][62] = 8'd23;
        rom[396][63] = 8'd3;
        rom[397][0] = -8'd43;
        rom[397][1] = -8'd1;
        rom[397][2] = -8'd46;
        rom[397][3] = 8'd27;
        rom[397][4] = 8'd1;
        rom[397][5] = 8'd2;
        rom[397][6] = 8'd0;
        rom[397][7] = 8'd24;
        rom[397][8] = -8'd3;
        rom[397][9] = -8'd2;
        rom[397][10] = -8'd11;
        rom[397][11] = -8'd23;
        rom[397][12] = -8'd22;
        rom[397][13] = -8'd7;
        rom[397][14] = -8'd57;
        rom[397][15] = 8'd5;
        rom[397][16] = -8'd6;
        rom[397][17] = 8'd15;
        rom[397][18] = -8'd6;
        rom[397][19] = 8'd3;
        rom[397][20] = 8'd1;
        rom[397][21] = -8'd17;
        rom[397][22] = -8'd23;
        rom[397][23] = 8'd10;
        rom[397][24] = -8'd5;
        rom[397][25] = 8'd29;
        rom[397][26] = 8'd11;
        rom[397][27] = 8'd25;
        rom[397][28] = 8'd3;
        rom[397][29] = -8'd8;
        rom[397][30] = -8'd50;
        rom[397][31] = 8'd1;
        rom[397][32] = -8'd7;
        rom[397][33] = 8'd9;
        rom[397][34] = -8'd39;
        rom[397][35] = -8'd26;
        rom[397][36] = 8'd3;
        rom[397][37] = 8'd22;
        rom[397][38] = -8'd41;
        rom[397][39] = -8'd2;
        rom[397][40] = 8'd18;
        rom[397][41] = -8'd1;
        rom[397][42] = -8'd13;
        rom[397][43] = 8'd25;
        rom[397][44] = -8'd7;
        rom[397][45] = 8'd11;
        rom[397][46] = -8'd18;
        rom[397][47] = -8'd12;
        rom[397][48] = -8'd48;
        rom[397][49] = -8'd13;
        rom[397][50] = -8'd42;
        rom[397][51] = -8'd53;
        rom[397][52] = 8'd31;
        rom[397][53] = -8'd7;
        rom[397][54] = 8'd4;
        rom[397][55] = 8'd10;
        rom[397][56] = -8'd30;
        rom[397][57] = -8'd5;
        rom[397][58] = -8'd2;
        rom[397][59] = -8'd16;
        rom[397][60] = 8'd20;
        rom[397][61] = -8'd28;
        rom[397][62] = -8'd10;
        rom[397][63] = -8'd29;
        rom[398][0] = -8'd19;
        rom[398][1] = 8'd16;
        rom[398][2] = -8'd20;
        rom[398][3] = -8'd13;
        rom[398][4] = 8'd13;
        rom[398][5] = -8'd24;
        rom[398][6] = -8'd27;
        rom[398][7] = -8'd50;
        rom[398][8] = 8'd35;
        rom[398][9] = -8'd35;
        rom[398][10] = 8'd31;
        rom[398][11] = 8'd17;
        rom[398][12] = 8'd7;
        rom[398][13] = -8'd14;
        rom[398][14] = 8'd2;
        rom[398][15] = -8'd23;
        rom[398][16] = -8'd105;
        rom[398][17] = -8'd32;
        rom[398][18] = 8'd12;
        rom[398][19] = 8'd31;
        rom[398][20] = -8'd3;
        rom[398][21] = 8'd36;
        rom[398][22] = 8'd13;
        rom[398][23] = -8'd5;
        rom[398][24] = -8'd5;
        rom[398][25] = 8'd59;
        rom[398][26] = 8'd29;
        rom[398][27] = -8'd20;
        rom[398][28] = -8'd9;
        rom[398][29] = 8'd17;
        rom[398][30] = -8'd20;
        rom[398][31] = 8'd12;
        rom[398][32] = 8'd21;
        rom[398][33] = -8'd31;
        rom[398][34] = 8'd34;
        rom[398][35] = -8'd26;
        rom[398][36] = 8'd3;
        rom[398][37] = 8'd12;
        rom[398][38] = 8'd48;
        rom[398][39] = -8'd5;
        rom[398][40] = -8'd1;
        rom[398][41] = 8'd21;
        rom[398][42] = -8'd9;
        rom[398][43] = -8'd11;
        rom[398][44] = 8'd11;
        rom[398][45] = 8'd9;
        rom[398][46] = -8'd27;
        rom[398][47] = -8'd41;
        rom[398][48] = -8'd1;
        rom[398][49] = 8'd20;
        rom[398][50] = -8'd3;
        rom[398][51] = 8'd27;
        rom[398][52] = 8'd5;
        rom[398][53] = 8'd30;
        rom[398][54] = 8'd13;
        rom[398][55] = 8'd7;
        rom[398][56] = 8'd7;
        rom[398][57] = 8'd5;
        rom[398][58] = -8'd6;
        rom[398][59] = -8'd36;
        rom[398][60] = -8'd5;
        rom[398][61] = -8'd1;
        rom[398][62] = 8'd17;
        rom[398][63] = 8'd11;
        rom[399][0] = 8'd3;
        rom[399][1] = 8'd5;
        rom[399][2] = 8'd11;
        rom[399][3] = -8'd16;
        rom[399][4] = 8'd3;
        rom[399][5] = -8'd9;
        rom[399][6] = -8'd16;
        rom[399][7] = -8'd19;
        rom[399][8] = 8'd12;
        rom[399][9] = -8'd34;
        rom[399][10] = -8'd28;
        rom[399][11] = -8'd11;
        rom[399][12] = 8'd14;
        rom[399][13] = -8'd16;
        rom[399][14] = 8'd1;
        rom[399][15] = 8'd3;
        rom[399][16] = -8'd30;
        rom[399][17] = 8'd3;
        rom[399][18] = 8'd15;
        rom[399][19] = -8'd5;
        rom[399][20] = -8'd13;
        rom[399][21] = -8'd28;
        rom[399][22] = -8'd6;
        rom[399][23] = 8'd7;
        rom[399][24] = -8'd25;
        rom[399][25] = -8'd37;
        rom[399][26] = 8'd10;
        rom[399][27] = -8'd21;
        rom[399][28] = -8'd35;
        rom[399][29] = 8'd14;
        rom[399][30] = -8'd8;
        rom[399][31] = -8'd38;
        rom[399][32] = 8'd28;
        rom[399][33] = 8'd0;
        rom[399][34] = 8'd9;
        rom[399][35] = 8'd21;
        rom[399][36] = 8'd11;
        rom[399][37] = -8'd25;
        rom[399][38] = 8'd10;
        rom[399][39] = 8'd24;
        rom[399][40] = -8'd8;
        rom[399][41] = 8'd9;
        rom[399][42] = 8'd5;
        rom[399][43] = 8'd1;
        rom[399][44] = 8'd18;
        rom[399][45] = 8'd8;
        rom[399][46] = -8'd7;
        rom[399][47] = 8'd0;
        rom[399][48] = 8'd9;
        rom[399][49] = 8'd10;
        rom[399][50] = -8'd15;
        rom[399][51] = 8'd41;
        rom[399][52] = 8'd3;
        rom[399][53] = 8'd18;
        rom[399][54] = 8'd5;
        rom[399][55] = -8'd47;
        rom[399][56] = -8'd27;
        rom[399][57] = -8'd13;
        rom[399][58] = -8'd4;
        rom[399][59] = -8'd32;
        rom[399][60] = 8'd10;
        rom[399][61] = -8'd70;
        rom[399][62] = 8'd1;
        rom[399][63] = -8'd24;
        rom[400][0] = 8'd2;
        rom[400][1] = 8'd9;
        rom[400][2] = -8'd8;
        rom[400][3] = 8'd0;
        rom[400][4] = -8'd1;
        rom[400][5] = -8'd1;
        rom[400][6] = -8'd8;
        rom[400][7] = -8'd9;
        rom[400][8] = 8'd3;
        rom[400][9] = 8'd9;
        rom[400][10] = -8'd3;
        rom[400][11] = 8'd0;
        rom[400][12] = 8'd4;
        rom[400][13] = 8'd6;
        rom[400][14] = -8'd1;
        rom[400][15] = -8'd4;
        rom[400][16] = 8'd3;
        rom[400][17] = -8'd2;
        rom[400][18] = 8'd5;
        rom[400][19] = -8'd4;
        rom[400][20] = 8'd5;
        rom[400][21] = -8'd4;
        rom[400][22] = -8'd6;
        rom[400][23] = -8'd1;
        rom[400][24] = 8'd6;
        rom[400][25] = -8'd4;
        rom[400][26] = -8'd8;
        rom[400][27] = -8'd8;
        rom[400][28] = 8'd3;
        rom[400][29] = -8'd7;
        rom[400][30] = -8'd5;
        rom[400][31] = 8'd0;
        rom[400][32] = -8'd8;
        rom[400][33] = -8'd8;
        rom[400][34] = 8'd1;
        rom[400][35] = 8'd3;
        rom[400][36] = 8'd1;
        rom[400][37] = 8'd8;
        rom[400][38] = -8'd3;
        rom[400][39] = 8'd8;
        rom[400][40] = -8'd9;
        rom[400][41] = 8'd7;
        rom[400][42] = -8'd4;
        rom[400][43] = 8'd4;
        rom[400][44] = 8'd1;
        rom[400][45] = 8'd5;
        rom[400][46] = -8'd1;
        rom[400][47] = 8'd5;
        rom[400][48] = 8'd7;
        rom[400][49] = 8'd3;
        rom[400][50] = -8'd6;
        rom[400][51] = 8'd6;
        rom[400][52] = -8'd3;
        rom[400][53] = 8'd2;
        rom[400][54] = -8'd5;
        rom[400][55] = 8'd4;
        rom[400][56] = 8'd1;
        rom[400][57] = 8'd0;
        rom[400][58] = 8'd10;
        rom[400][59] = 8'd4;
        rom[400][60] = -8'd4;
        rom[400][61] = -8'd9;
        rom[400][62] = 8'd8;
        rom[400][63] = -8'd3;
        rom[401][0] = 8'd20;
        rom[401][1] = 8'd21;
        rom[401][2] = 8'd11;
        rom[401][3] = -8'd10;
        rom[401][4] = 8'd37;
        rom[401][5] = 8'd18;
        rom[401][6] = 8'd14;
        rom[401][7] = -8'd42;
        rom[401][8] = -8'd18;
        rom[401][9] = 8'd0;
        rom[401][10] = 8'd17;
        rom[401][11] = -8'd20;
        rom[401][12] = -8'd32;
        rom[401][13] = -8'd16;
        rom[401][14] = 8'd38;
        rom[401][15] = 8'd5;
        rom[401][16] = -8'd13;
        rom[401][17] = -8'd38;
        rom[401][18] = -8'd28;
        rom[401][19] = -8'd29;
        rom[401][20] = -8'd6;
        rom[401][21] = -8'd18;
        rom[401][22] = -8'd3;
        rom[401][23] = -8'd6;
        rom[401][24] = 8'd4;
        rom[401][25] = -8'd42;
        rom[401][26] = -8'd11;
        rom[401][27] = -8'd15;
        rom[401][28] = -8'd38;
        rom[401][29] = 8'd37;
        rom[401][30] = -8'd8;
        rom[401][31] = 8'd24;
        rom[401][32] = 8'd21;
        rom[401][33] = 8'd21;
        rom[401][34] = -8'd34;
        rom[401][35] = -8'd11;
        rom[401][36] = -8'd85;
        rom[401][37] = 8'd26;
        rom[401][38] = -8'd48;
        rom[401][39] = 8'd3;
        rom[401][40] = 8'd18;
        rom[401][41] = -8'd27;
        rom[401][42] = 8'd3;
        rom[401][43] = 8'd16;
        rom[401][44] = 8'd6;
        rom[401][45] = 8'd45;
        rom[401][46] = 8'd30;
        rom[401][47] = 8'd26;
        rom[401][48] = 8'd9;
        rom[401][49] = -8'd10;
        rom[401][50] = 8'd2;
        rom[401][51] = 8'd4;
        rom[401][52] = 8'd38;
        rom[401][53] = -8'd5;
        rom[401][54] = -8'd19;
        rom[401][55] = -8'd2;
        rom[401][56] = -8'd7;
        rom[401][57] = 8'd46;
        rom[401][58] = -8'd41;
        rom[401][59] = 8'd31;
        rom[401][60] = 8'd15;
        rom[401][61] = -8'd11;
        rom[401][62] = 8'd7;
        rom[401][63] = -8'd4;
        rom[402][0] = 8'd26;
        rom[402][1] = -8'd30;
        rom[402][2] = 8'd0;
        rom[402][3] = -8'd34;
        rom[402][4] = 8'd9;
        rom[402][5] = -8'd33;
        rom[402][6] = 8'd20;
        rom[402][7] = -8'd56;
        rom[402][8] = 8'd13;
        rom[402][9] = -8'd12;
        rom[402][10] = 8'd10;
        rom[402][11] = 8'd1;
        rom[402][12] = -8'd13;
        rom[402][13] = -8'd48;
        rom[402][14] = 8'd16;
        rom[402][15] = -8'd18;
        rom[402][16] = -8'd109;
        rom[402][17] = -8'd37;
        rom[402][18] = -8'd21;
        rom[402][19] = 8'd10;
        rom[402][20] = -8'd7;
        rom[402][21] = 8'd14;
        rom[402][22] = -8'd15;
        rom[402][23] = 8'd2;
        rom[402][24] = -8'd5;
        rom[402][25] = -8'd18;
        rom[402][26] = -8'd69;
        rom[402][27] = -8'd7;
        rom[402][28] = 8'd15;
        rom[402][29] = -8'd66;
        rom[402][30] = -8'd35;
        rom[402][31] = -8'd14;
        rom[402][32] = 8'd14;
        rom[402][33] = -8'd39;
        rom[402][34] = -8'd14;
        rom[402][35] = 8'd7;
        rom[402][36] = -8'd16;
        rom[402][37] = -8'd32;
        rom[402][38] = -8'd40;
        rom[402][39] = 8'd43;
        rom[402][40] = -8'd29;
        rom[402][41] = 8'd6;
        rom[402][42] = 8'd0;
        rom[402][43] = 8'd4;
        rom[402][44] = 8'd6;
        rom[402][45] = -8'd91;
        rom[402][46] = -8'd2;
        rom[402][47] = -8'd13;
        rom[402][48] = -8'd12;
        rom[402][49] = -8'd44;
        rom[402][50] = -8'd13;
        rom[402][51] = -8'd4;
        rom[402][52] = -8'd26;
        rom[402][53] = 8'd6;
        rom[402][54] = -8'd11;
        rom[402][55] = 8'd33;
        rom[402][56] = -8'd13;
        rom[402][57] = -8'd14;
        rom[402][58] = -8'd26;
        rom[402][59] = -8'd19;
        rom[402][60] = -8'd39;
        rom[402][61] = 8'd36;
        rom[402][62] = -8'd3;
        rom[402][63] = 8'd30;
        rom[403][0] = -8'd1;
        rom[403][1] = -8'd7;
        rom[403][2] = 8'd22;
        rom[403][3] = -8'd45;
        rom[403][4] = -8'd13;
        rom[403][5] = 8'd4;
        rom[403][6] = -8'd15;
        rom[403][7] = 8'd37;
        rom[403][8] = -8'd60;
        rom[403][9] = -8'd16;
        rom[403][10] = 8'd4;
        rom[403][11] = -8'd35;
        rom[403][12] = -8'd12;
        rom[403][13] = 8'd17;
        rom[403][14] = -8'd33;
        rom[403][15] = 8'd45;
        rom[403][16] = 8'd30;
        rom[403][17] = -8'd29;
        rom[403][18] = 8'd6;
        rom[403][19] = -8'd20;
        rom[403][20] = -8'd4;
        rom[403][21] = -8'd9;
        rom[403][22] = -8'd5;
        rom[403][23] = 8'd9;
        rom[403][24] = -8'd21;
        rom[403][25] = 8'd16;
        rom[403][26] = -8'd38;
        rom[403][27] = -8'd30;
        rom[403][28] = -8'd5;
        rom[403][29] = 8'd5;
        rom[403][30] = 8'd27;
        rom[403][31] = -8'd47;
        rom[403][32] = 8'd21;
        rom[403][33] = 8'd4;
        rom[403][34] = 8'd9;
        rom[403][35] = -8'd7;
        rom[403][36] = 8'd0;
        rom[403][37] = -8'd53;
        rom[403][38] = -8'd35;
        rom[403][39] = 8'd34;
        rom[403][40] = 8'd12;
        rom[403][41] = -8'd24;
        rom[403][42] = 8'd16;
        rom[403][43] = 8'd21;
        rom[403][44] = 8'd36;
        rom[403][45] = 8'd5;
        rom[403][46] = 8'd12;
        rom[403][47] = 8'd38;
        rom[403][48] = -8'd31;
        rom[403][49] = -8'd18;
        rom[403][50] = 8'd2;
        rom[403][51] = 8'd14;
        rom[403][52] = 8'd31;
        rom[403][53] = 8'd9;
        rom[403][54] = -8'd40;
        rom[403][55] = -8'd38;
        rom[403][56] = -8'd13;
        rom[403][57] = 8'd25;
        rom[403][58] = -8'd23;
        rom[403][59] = -8'd5;
        rom[403][60] = 8'd10;
        rom[403][61] = -8'd18;
        rom[403][62] = 8'd9;
        rom[403][63] = 8'd3;
        rom[404][0] = 8'd2;
        rom[404][1] = -8'd21;
        rom[404][2] = -8'd63;
        rom[404][3] = 8'd11;
        rom[404][4] = -8'd47;
        rom[404][5] = 8'd2;
        rom[404][6] = 8'd13;
        rom[404][7] = 8'd20;
        rom[404][8] = -8'd40;
        rom[404][9] = -8'd45;
        rom[404][10] = -8'd20;
        rom[404][11] = 8'd19;
        rom[404][12] = 8'd7;
        rom[404][13] = -8'd51;
        rom[404][14] = -8'd30;
        rom[404][15] = -8'd31;
        rom[404][16] = -8'd68;
        rom[404][17] = -8'd29;
        rom[404][18] = -8'd30;
        rom[404][19] = -8'd24;
        rom[404][20] = -8'd8;
        rom[404][21] = 8'd28;
        rom[404][22] = -8'd11;
        rom[404][23] = -8'd12;
        rom[404][24] = 8'd8;
        rom[404][25] = -8'd2;
        rom[404][26] = 8'd24;
        rom[404][27] = 8'd1;
        rom[404][28] = -8'd24;
        rom[404][29] = -8'd86;
        rom[404][30] = -8'd30;
        rom[404][31] = -8'd39;
        rom[404][32] = -8'd13;
        rom[404][33] = -8'd38;
        rom[404][34] = 8'd38;
        rom[404][35] = 8'd5;
        rom[404][36] = -8'd38;
        rom[404][37] = -8'd75;
        rom[404][38] = 8'd21;
        rom[404][39] = 8'd27;
        rom[404][40] = 8'd14;
        rom[404][41] = -8'd21;
        rom[404][42] = -8'd23;
        rom[404][43] = -8'd2;
        rom[404][44] = -8'd11;
        rom[404][45] = -8'd38;
        rom[404][46] = 8'd12;
        rom[404][47] = -8'd8;
        rom[404][48] = -8'd36;
        rom[404][49] = 8'd9;
        rom[404][50] = -8'd110;
        rom[404][51] = 8'd34;
        rom[404][52] = 8'd19;
        rom[404][53] = -8'd12;
        rom[404][54] = 8'd35;
        rom[404][55] = -8'd28;
        rom[404][56] = -8'd4;
        rom[404][57] = -8'd12;
        rom[404][58] = 8'd3;
        rom[404][59] = -8'd15;
        rom[404][60] = -8'd11;
        rom[404][61] = -8'd8;
        rom[404][62] = -8'd8;
        rom[404][63] = -8'd20;
        rom[405][0] = 8'd6;
        rom[405][1] = 8'd3;
        rom[405][2] = 8'd4;
        rom[405][3] = 8'd1;
        rom[405][4] = -8'd8;
        rom[405][5] = 8'd6;
        rom[405][6] = -8'd8;
        rom[405][7] = -8'd7;
        rom[405][8] = -8'd5;
        rom[405][9] = 8'd8;
        rom[405][10] = 8'd1;
        rom[405][11] = 8'd6;
        rom[405][12] = 8'd3;
        rom[405][13] = -8'd6;
        rom[405][14] = -8'd1;
        rom[405][15] = 8'd6;
        rom[405][16] = 8'd6;
        rom[405][17] = 8'd5;
        rom[405][18] = 8'd7;
        rom[405][19] = 8'd5;
        rom[405][20] = 8'd4;
        rom[405][21] = -8'd1;
        rom[405][22] = -8'd3;
        rom[405][23] = 8'd0;
        rom[405][24] = 8'd8;
        rom[405][25] = 8'd7;
        rom[405][26] = -8'd1;
        rom[405][27] = 8'd4;
        rom[405][28] = 8'd6;
        rom[405][29] = -8'd2;
        rom[405][30] = 8'd1;
        rom[405][31] = 8'd0;
        rom[405][32] = 8'd4;
        rom[405][33] = 8'd3;
        rom[405][34] = -8'd11;
        rom[405][35] = 8'd0;
        rom[405][36] = 8'd0;
        rom[405][37] = 8'd6;
        rom[405][38] = 8'd4;
        rom[405][39] = -8'd1;
        rom[405][40] = -8'd7;
        rom[405][41] = 8'd3;
        rom[405][42] = 8'd2;
        rom[405][43] = 8'd0;
        rom[405][44] = 8'd3;
        rom[405][45] = -8'd3;
        rom[405][46] = -8'd6;
        rom[405][47] = 8'd2;
        rom[405][48] = -8'd8;
        rom[405][49] = 8'd6;
        rom[405][50] = -8'd7;
        rom[405][51] = -8'd7;
        rom[405][52] = 8'd3;
        rom[405][53] = 8'd5;
        rom[405][54] = -8'd3;
        rom[405][55] = 8'd0;
        rom[405][56] = 8'd6;
        rom[405][57] = 8'd1;
        rom[405][58] = 8'd2;
        rom[405][59] = -8'd5;
        rom[405][60] = 8'd1;
        rom[405][61] = 8'd1;
        rom[405][62] = 8'd4;
        rom[405][63] = 8'd3;
        rom[406][0] = -8'd78;
        rom[406][1] = -8'd2;
        rom[406][2] = -8'd20;
        rom[406][3] = 8'd22;
        rom[406][4] = 8'd3;
        rom[406][5] = 8'd5;
        rom[406][6] = -8'd12;
        rom[406][7] = -8'd29;
        rom[406][8] = 8'd11;
        rom[406][9] = -8'd2;
        rom[406][10] = 8'd5;
        rom[406][11] = -8'd46;
        rom[406][12] = -8'd13;
        rom[406][13] = 8'd27;
        rom[406][14] = 8'd33;
        rom[406][15] = 8'd1;
        rom[406][16] = -8'd3;
        rom[406][17] = 8'd4;
        rom[406][18] = -8'd40;
        rom[406][19] = 8'd21;
        rom[406][20] = -8'd1;
        rom[406][21] = -8'd24;
        rom[406][22] = -8'd17;
        rom[406][23] = 8'd22;
        rom[406][24] = -8'd16;
        rom[406][25] = -8'd10;
        rom[406][26] = 8'd4;
        rom[406][27] = 8'd2;
        rom[406][28] = 8'd17;
        rom[406][29] = -8'd1;
        rom[406][30] = -8'd5;
        rom[406][31] = 8'd9;
        rom[406][32] = 8'd16;
        rom[406][33] = -8'd6;
        rom[406][34] = -8'd2;
        rom[406][35] = 8'd12;
        rom[406][36] = -8'd36;
        rom[406][37] = -8'd3;
        rom[406][38] = -8'd27;
        rom[406][39] = 8'd19;
        rom[406][40] = 8'd16;
        rom[406][41] = 8'd28;
        rom[406][42] = -8'd32;
        rom[406][43] = 8'd3;
        rom[406][44] = -8'd31;
        rom[406][45] = -8'd52;
        rom[406][46] = 8'd18;
        rom[406][47] = -8'd25;
        rom[406][48] = -8'd10;
        rom[406][49] = -8'd3;
        rom[406][50] = -8'd12;
        rom[406][51] = -8'd13;
        rom[406][52] = -8'd5;
        rom[406][53] = 8'd36;
        rom[406][54] = -8'd11;
        rom[406][55] = -8'd19;
        rom[406][56] = 8'd7;
        rom[406][57] = 8'd3;
        rom[406][58] = 8'd22;
        rom[406][59] = -8'd5;
        rom[406][60] = -8'd6;
        rom[406][61] = 8'd8;
        rom[406][62] = 8'd14;
        rom[406][63] = -8'd10;
        rom[407][0] = 8'd2;
        rom[407][1] = -8'd4;
        rom[407][2] = 8'd0;
        rom[407][3] = 8'd5;
        rom[407][4] = -8'd6;
        rom[407][5] = -8'd5;
        rom[407][6] = 8'd7;
        rom[407][7] = 8'd10;
        rom[407][8] = -8'd5;
        rom[407][9] = 8'd11;
        rom[407][10] = -8'd19;
        rom[407][11] = -8'd16;
        rom[407][12] = 8'd22;
        rom[407][13] = 8'd41;
        rom[407][14] = -8'd14;
        rom[407][15] = -8'd10;
        rom[407][16] = -8'd24;
        rom[407][17] = 8'd11;
        rom[407][18] = 8'd40;
        rom[407][19] = -8'd6;
        rom[407][20] = -8'd2;
        rom[407][21] = -8'd7;
        rom[407][22] = 8'd20;
        rom[407][23] = -8'd31;
        rom[407][24] = -8'd13;
        rom[407][25] = -8'd4;
        rom[407][26] = -8'd23;
        rom[407][27] = -8'd6;
        rom[407][28] = -8'd8;
        rom[407][29] = -8'd20;
        rom[407][30] = 8'd46;
        rom[407][31] = -8'd2;
        rom[407][32] = 8'd24;
        rom[407][33] = -8'd46;
        rom[407][34] = 8'd20;
        rom[407][35] = 8'd42;
        rom[407][36] = -8'd40;
        rom[407][37] = -8'd36;
        rom[407][38] = 8'd3;
        rom[407][39] = -8'd1;
        rom[407][40] = -8'd15;
        rom[407][41] = -8'd12;
        rom[407][42] = -8'd5;
        rom[407][43] = 8'd16;
        rom[407][44] = -8'd23;
        rom[407][45] = -8'd13;
        rom[407][46] = -8'd12;
        rom[407][47] = 8'd21;
        rom[407][48] = 8'd20;
        rom[407][49] = 8'd21;
        rom[407][50] = -8'd14;
        rom[407][51] = -8'd8;
        rom[407][52] = -8'd17;
        rom[407][53] = -8'd1;
        rom[407][54] = -8'd28;
        rom[407][55] = 8'd33;
        rom[407][56] = -8'd8;
        rom[407][57] = 8'd3;
        rom[407][58] = -8'd28;
        rom[407][59] = -8'd8;
        rom[407][60] = -8'd20;
        rom[407][61] = 8'd0;
        rom[407][62] = -8'd19;
        rom[407][63] = 8'd18;
        rom[408][0] = -8'd27;
        rom[408][1] = -8'd5;
        rom[408][2] = 8'd4;
        rom[408][3] = 8'd16;
        rom[408][4] = 8'd65;
        rom[408][5] = -8'd4;
        rom[408][6] = 8'd38;
        rom[408][7] = 8'd27;
        rom[408][8] = -8'd35;
        rom[408][9] = 8'd34;
        rom[408][10] = 8'd35;
        rom[408][11] = 8'd17;
        rom[408][12] = 8'd11;
        rom[408][13] = 8'd10;
        rom[408][14] = 8'd10;
        rom[408][15] = -8'd6;
        rom[408][16] = 8'd4;
        rom[408][17] = -8'd15;
        rom[408][18] = 8'd23;
        rom[408][19] = 8'd30;
        rom[408][20] = -8'd6;
        rom[408][21] = -8'd20;
        rom[408][22] = 8'd36;
        rom[408][23] = 8'd13;
        rom[408][24] = 8'd0;
        rom[408][25] = -8'd34;
        rom[408][26] = 8'd31;
        rom[408][27] = -8'd26;
        rom[408][28] = 8'd34;
        rom[408][29] = -8'd41;
        rom[408][30] = 8'd26;
        rom[408][31] = -8'd25;
        rom[408][32] = 8'd41;
        rom[408][33] = -8'd9;
        rom[408][34] = -8'd18;
        rom[408][35] = 8'd39;
        rom[408][36] = -8'd30;
        rom[408][37] = 8'd3;
        rom[408][38] = -8'd7;
        rom[408][39] = 8'd30;
        rom[408][40] = 8'd14;
        rom[408][41] = 8'd7;
        rom[408][42] = 8'd18;
        rom[408][43] = -8'd3;
        rom[408][44] = -8'd57;
        rom[408][45] = -8'd6;
        rom[408][46] = 8'd38;
        rom[408][47] = 8'd36;
        rom[408][48] = 8'd36;
        rom[408][49] = -8'd13;
        rom[408][50] = 8'd6;
        rom[408][51] = -8'd22;
        rom[408][52] = 8'd12;
        rom[408][53] = 8'd23;
        rom[408][54] = 8'd29;
        rom[408][55] = -8'd15;
        rom[408][56] = 8'd1;
        rom[408][57] = 8'd28;
        rom[408][58] = -8'd59;
        rom[408][59] = 8'd4;
        rom[408][60] = -8'd4;
        rom[408][61] = 8'd38;
        rom[408][62] = -8'd15;
        rom[408][63] = -8'd2;
        rom[409][0] = 8'd11;
        rom[409][1] = -8'd19;
        rom[409][2] = 8'd16;
        rom[409][3] = -8'd7;
        rom[409][4] = -8'd14;
        rom[409][5] = -8'd1;
        rom[409][6] = 8'd21;
        rom[409][7] = 8'd19;
        rom[409][8] = 8'd8;
        rom[409][9] = 8'd12;
        rom[409][10] = 8'd8;
        rom[409][11] = -8'd2;
        rom[409][12] = 8'd3;
        rom[409][13] = -8'd33;
        rom[409][14] = 8'd47;
        rom[409][15] = 8'd16;
        rom[409][16] = -8'd10;
        rom[409][17] = 8'd20;
        rom[409][18] = -8'd42;
        rom[409][19] = 8'd9;
        rom[409][20] = -8'd8;
        rom[409][21] = 8'd3;
        rom[409][22] = 8'd25;
        rom[409][23] = 8'd7;
        rom[409][24] = 8'd25;
        rom[409][25] = 8'd7;
        rom[409][26] = 8'd9;
        rom[409][27] = -8'd21;
        rom[409][28] = -8'd13;
        rom[409][29] = 8'd0;
        rom[409][30] = -8'd12;
        rom[409][31] = 8'd10;
        rom[409][32] = 8'd14;
        rom[409][33] = -8'd24;
        rom[409][34] = 8'd1;
        rom[409][35] = -8'd4;
        rom[409][36] = 8'd18;
        rom[409][37] = 8'd11;
        rom[409][38] = -8'd39;
        rom[409][39] = -8'd21;
        rom[409][40] = -8'd30;
        rom[409][41] = -8'd15;
        rom[409][42] = 8'd41;
        rom[409][43] = -8'd9;
        rom[409][44] = 8'd11;
        rom[409][45] = -8'd39;
        rom[409][46] = 8'd3;
        rom[409][47] = 8'd18;
        rom[409][48] = -8'd52;
        rom[409][49] = -8'd26;
        rom[409][50] = 8'd17;
        rom[409][51] = 8'd8;
        rom[409][52] = -8'd8;
        rom[409][53] = -8'd28;
        rom[409][54] = 8'd9;
        rom[409][55] = 8'd29;
        rom[409][56] = -8'd24;
        rom[409][57] = 8'd45;
        rom[409][58] = -8'd1;
        rom[409][59] = -8'd5;
        rom[409][60] = 8'd56;
        rom[409][61] = -8'd26;
        rom[409][62] = 8'd1;
        rom[409][63] = 8'd32;
        rom[410][0] = 8'd39;
        rom[410][1] = -8'd33;
        rom[410][2] = -8'd9;
        rom[410][3] = 8'd2;
        rom[410][4] = -8'd2;
        rom[410][5] = 8'd0;
        rom[410][6] = 8'd3;
        rom[410][7] = -8'd4;
        rom[410][8] = 8'd2;
        rom[410][9] = 8'd37;
        rom[410][10] = 8'd38;
        rom[410][11] = 8'd22;
        rom[410][12] = -8'd38;
        rom[410][13] = -8'd37;
        rom[410][14] = 8'd8;
        rom[410][15] = -8'd2;
        rom[410][16] = 8'd3;
        rom[410][17] = 8'd44;
        rom[410][18] = 8'd44;
        rom[410][19] = -8'd23;
        rom[410][20] = -8'd1;
        rom[410][21] = -8'd13;
        rom[410][22] = 8'd0;
        rom[410][23] = -8'd10;
        rom[410][24] = -8'd35;
        rom[410][25] = -8'd13;
        rom[410][26] = -8'd21;
        rom[410][27] = -8'd86;
        rom[410][28] = -8'd33;
        rom[410][29] = -8'd34;
        rom[410][30] = 8'd30;
        rom[410][31] = 8'd3;
        rom[410][32] = 8'd11;
        rom[410][33] = -8'd8;
        rom[410][34] = 8'd47;
        rom[410][35] = -8'd54;
        rom[410][36] = 8'd8;
        rom[410][37] = 8'd7;
        rom[410][38] = 8'd36;
        rom[410][39] = 8'd10;
        rom[410][40] = 8'd1;
        rom[410][41] = -8'd11;
        rom[410][42] = -8'd30;
        rom[410][43] = -8'd26;
        rom[410][44] = 8'd11;
        rom[410][45] = 8'd14;
        rom[410][46] = -8'd112;
        rom[410][47] = -8'd15;
        rom[410][48] = 8'd43;
        rom[410][49] = -8'd26;
        rom[410][50] = -8'd53;
        rom[410][51] = 8'd8;
        rom[410][52] = 8'd14;
        rom[410][53] = 8'd37;
        rom[410][54] = 8'd11;
        rom[410][55] = 8'd44;
        rom[410][56] = 8'd13;
        rom[410][57] = 8'd50;
        rom[410][58] = -8'd55;
        rom[410][59] = 8'd22;
        rom[410][60] = 8'd32;
        rom[410][61] = 8'd3;
        rom[410][62] = 8'd4;
        rom[410][63] = 8'd0;
        rom[411][0] = 8'd6;
        rom[411][1] = 8'd72;
        rom[411][2] = 8'd52;
        rom[411][3] = -8'd1;
        rom[411][4] = 8'd4;
        rom[411][5] = 8'd41;
        rom[411][6] = 8'd8;
        rom[411][7] = 8'd0;
        rom[411][8] = 8'd15;
        rom[411][9] = 8'd20;
        rom[411][10] = -8'd3;
        rom[411][11] = 8'd38;
        rom[411][12] = -8'd28;
        rom[411][13] = -8'd5;
        rom[411][14] = 8'd9;
        rom[411][15] = 8'd12;
        rom[411][16] = -8'd10;
        rom[411][17] = -8'd8;
        rom[411][18] = 8'd8;
        rom[411][19] = 8'd29;
        rom[411][20] = -8'd5;
        rom[411][21] = -8'd20;
        rom[411][22] = -8'd23;
        rom[411][23] = 8'd17;
        rom[411][24] = 8'd26;
        rom[411][25] = 8'd38;
        rom[411][26] = -8'd5;
        rom[411][27] = -8'd18;
        rom[411][28] = 8'd10;
        rom[411][29] = 8'd44;
        rom[411][30] = -8'd38;
        rom[411][31] = 8'd36;
        rom[411][32] = -8'd4;
        rom[411][33] = 8'd18;
        rom[411][34] = -8'd11;
        rom[411][35] = -8'd1;
        rom[411][36] = 8'd0;
        rom[411][37] = -8'd28;
        rom[411][38] = -8'd2;
        rom[411][39] = -8'd6;
        rom[411][40] = -8'd32;
        rom[411][41] = 8'd12;
        rom[411][42] = 8'd29;
        rom[411][43] = -8'd3;
        rom[411][44] = 8'd12;
        rom[411][45] = -8'd15;
        rom[411][46] = 8'd44;
        rom[411][47] = -8'd50;
        rom[411][48] = 8'd18;
        rom[411][49] = -8'd13;
        rom[411][50] = 8'd15;
        rom[411][51] = -8'd1;
        rom[411][52] = 8'd26;
        rom[411][53] = 8'd4;
        rom[411][54] = -8'd10;
        rom[411][55] = -8'd27;
        rom[411][56] = -8'd10;
        rom[411][57] = 8'd26;
        rom[411][58] = 8'd16;
        rom[411][59] = -8'd6;
        rom[411][60] = -8'd16;
        rom[411][61] = 8'd28;
        rom[411][62] = -8'd3;
        rom[411][63] = -8'd7;
        rom[412][0] = -8'd32;
        rom[412][1] = -8'd19;
        rom[412][2] = 8'd39;
        rom[412][3] = 8'd20;
        rom[412][4] = -8'd11;
        rom[412][5] = -8'd53;
        rom[412][6] = 8'd7;
        rom[412][7] = 8'd21;
        rom[412][8] = -8'd1;
        rom[412][9] = -8'd4;
        rom[412][10] = 8'd12;
        rom[412][11] = 8'd18;
        rom[412][12] = 8'd9;
        rom[412][13] = 8'd8;
        rom[412][14] = 8'd8;
        rom[412][15] = 8'd12;
        rom[412][16] = 8'd13;
        rom[412][17] = 8'd2;
        rom[412][18] = -8'd19;
        rom[412][19] = -8'd20;
        rom[412][20] = -8'd10;
        rom[412][21] = 8'd14;
        rom[412][22] = 8'd8;
        rom[412][23] = -8'd11;
        rom[412][24] = -8'd27;
        rom[412][25] = 8'd34;
        rom[412][26] = -8'd34;
        rom[412][27] = 8'd19;
        rom[412][28] = -8'd7;
        rom[412][29] = -8'd15;
        rom[412][30] = -8'd10;
        rom[412][31] = -8'd14;
        rom[412][32] = -8'd28;
        rom[412][33] = -8'd43;
        rom[412][34] = -8'd12;
        rom[412][35] = -8'd48;
        rom[412][36] = -8'd8;
        rom[412][37] = -8'd46;
        rom[412][38] = -8'd29;
        rom[412][39] = 8'd16;
        rom[412][40] = -8'd20;
        rom[412][41] = -8'd66;
        rom[412][42] = 8'd7;
        rom[412][43] = 8'd26;
        rom[412][44] = 8'd21;
        rom[412][45] = 8'd31;
        rom[412][46] = -8'd2;
        rom[412][47] = 8'd8;
        rom[412][48] = 8'd31;
        rom[412][49] = 8'd14;
        rom[412][50] = 8'd41;
        rom[412][51] = 8'd22;
        rom[412][52] = 8'd15;
        rom[412][53] = 8'd21;
        rom[412][54] = 8'd10;
        rom[412][55] = 8'd8;
        rom[412][56] = 8'd38;
        rom[412][57] = -8'd17;
        rom[412][58] = -8'd51;
        rom[412][59] = -8'd5;
        rom[412][60] = -8'd67;
        rom[412][61] = -8'd19;
        rom[412][62] = 8'd2;
        rom[412][63] = 8'd12;
        rom[413][0] = 8'd58;
        rom[413][1] = -8'd6;
        rom[413][2] = -8'd14;
        rom[413][3] = 8'd14;
        rom[413][4] = -8'd47;
        rom[413][5] = -8'd13;
        rom[413][6] = -8'd40;
        rom[413][7] = 8'd23;
        rom[413][8] = 8'd0;
        rom[413][9] = -8'd16;
        rom[413][10] = 8'd83;
        rom[413][11] = -8'd21;
        rom[413][12] = 8'd16;
        rom[413][13] = 8'd1;
        rom[413][14] = -8'd47;
        rom[413][15] = 8'd14;
        rom[413][16] = 8'd16;
        rom[413][17] = 8'd2;
        rom[413][18] = -8'd14;
        rom[413][19] = -8'd3;
        rom[413][20] = -8'd2;
        rom[413][21] = 8'd20;
        rom[413][22] = 8'd33;
        rom[413][23] = 8'd29;
        rom[413][24] = -8'd8;
        rom[413][25] = -8'd13;
        rom[413][26] = -8'd42;
        rom[413][27] = -8'd50;
        rom[413][28] = -8'd6;
        rom[413][29] = 8'd6;
        rom[413][30] = -8'd7;
        rom[413][31] = 8'd0;
        rom[413][32] = 8'd18;
        rom[413][33] = 8'd36;
        rom[413][34] = 8'd5;
        rom[413][35] = 8'd17;
        rom[413][36] = -8'd8;
        rom[413][37] = -8'd33;
        rom[413][38] = -8'd41;
        rom[413][39] = -8'd17;
        rom[413][40] = -8'd15;
        rom[413][41] = -8'd19;
        rom[413][42] = -8'd32;
        rom[413][43] = -8'd34;
        rom[413][44] = -8'd20;
        rom[413][45] = -8'd13;
        rom[413][46] = 8'd15;
        rom[413][47] = 8'd5;
        rom[413][48] = 8'd6;
        rom[413][49] = 8'd21;
        rom[413][50] = 8'd8;
        rom[413][51] = 8'd59;
        rom[413][52] = 8'd21;
        rom[413][53] = 8'd1;
        rom[413][54] = -8'd13;
        rom[413][55] = -8'd23;
        rom[413][56] = -8'd8;
        rom[413][57] = 8'd8;
        rom[413][58] = -8'd17;
        rom[413][59] = -8'd2;
        rom[413][60] = -8'd18;
        rom[413][61] = -8'd12;
        rom[413][62] = -8'd1;
        rom[413][63] = 8'd23;
        rom[414][0] = -8'd15;
        rom[414][1] = -8'd15;
        rom[414][2] = -8'd36;
        rom[414][3] = -8'd5;
        rom[414][4] = 8'd9;
        rom[414][5] = -8'd26;
        rom[414][6] = -8'd6;
        rom[414][7] = -8'd73;
        rom[414][8] = 8'd21;
        rom[414][9] = 8'd0;
        rom[414][10] = 8'd17;
        rom[414][11] = -8'd16;
        rom[414][12] = 8'd4;
        rom[414][13] = -8'd4;
        rom[414][14] = -8'd63;
        rom[414][15] = -8'd38;
        rom[414][16] = 8'd18;
        rom[414][17] = -8'd37;
        rom[414][18] = -8'd34;
        rom[414][19] = -8'd15;
        rom[414][20] = -8'd6;
        rom[414][21] = -8'd1;
        rom[414][22] = 8'd5;
        rom[414][23] = -8'd6;
        rom[414][24] = -8'd17;
        rom[414][25] = -8'd29;
        rom[414][26] = 8'd22;
        rom[414][27] = -8'd4;
        rom[414][28] = 8'd6;
        rom[414][29] = -8'd52;
        rom[414][30] = 8'd1;
        rom[414][31] = -8'd30;
        rom[414][32] = 8'd1;
        rom[414][33] = -8'd32;
        rom[414][34] = -8'd37;
        rom[414][35] = 8'd9;
        rom[414][36] = -8'd12;
        rom[414][37] = 8'd4;
        rom[414][38] = -8'd21;
        rom[414][39] = 8'd33;
        rom[414][40] = 8'd11;
        rom[414][41] = 8'd9;
        rom[414][42] = -8'd40;
        rom[414][43] = 8'd45;
        rom[414][44] = -8'd12;
        rom[414][45] = -8'd28;
        rom[414][46] = -8'd8;
        rom[414][47] = 8'd11;
        rom[414][48] = -8'd15;
        rom[414][49] = 8'd6;
        rom[414][50] = -8'd27;
        rom[414][51] = -8'd54;
        rom[414][52] = 8'd6;
        rom[414][53] = -8'd63;
        rom[414][54] = -8'd13;
        rom[414][55] = 8'd40;
        rom[414][56] = -8'd13;
        rom[414][57] = -8'd5;
        rom[414][58] = -8'd11;
        rom[414][59] = 8'd27;
        rom[414][60] = 8'd5;
        rom[414][61] = 8'd9;
        rom[414][62] = 8'd13;
        rom[414][63] = -8'd17;
        rom[415][0] = 8'd39;
        rom[415][1] = -8'd12;
        rom[415][2] = 8'd31;
        rom[415][3] = 8'd27;
        rom[415][4] = -8'd75;
        rom[415][5] = -8'd46;
        rom[415][6] = -8'd61;
        rom[415][7] = -8'd19;
        rom[415][8] = 8'd8;
        rom[415][9] = -8'd13;
        rom[415][10] = 8'd48;
        rom[415][11] = 8'd6;
        rom[415][12] = 8'd5;
        rom[415][13] = -8'd39;
        rom[415][14] = -8'd3;
        rom[415][15] = 8'd39;
        rom[415][16] = -8'd42;
        rom[415][17] = -8'd8;
        rom[415][18] = -8'd1;
        rom[415][19] = -8'd31;
        rom[415][20] = -8'd9;
        rom[415][21] = -8'd2;
        rom[415][22] = -8'd23;
        rom[415][23] = -8'd4;
        rom[415][24] = -8'd23;
        rom[415][25] = -8'd21;
        rom[415][26] = 8'd13;
        rom[415][27] = -8'd54;
        rom[415][28] = -8'd3;
        rom[415][29] = 8'd23;
        rom[415][30] = 8'd8;
        rom[415][31] = 8'd16;
        rom[415][32] = 8'd27;
        rom[415][33] = 8'd12;
        rom[415][34] = 8'd11;
        rom[415][35] = -8'd19;
        rom[415][36] = -8'd14;
        rom[415][37] = -8'd13;
        rom[415][38] = 8'd9;
        rom[415][39] = -8'd28;
        rom[415][40] = 8'd1;
        rom[415][41] = -8'd14;
        rom[415][42] = 8'd4;
        rom[415][43] = -8'd29;
        rom[415][44] = 8'd16;
        rom[415][45] = -8'd41;
        rom[415][46] = -8'd10;
        rom[415][47] = -8'd13;
        rom[415][48] = -8'd50;
        rom[415][49] = -8'd12;
        rom[415][50] = -8'd13;
        rom[415][51] = -8'd32;
        rom[415][52] = 8'd19;
        rom[415][53] = 8'd23;
        rom[415][54] = -8'd8;
        rom[415][55] = 8'd26;
        rom[415][56] = 8'd60;
        rom[415][57] = 8'd5;
        rom[415][58] = 8'd47;
        rom[415][59] = 8'd25;
        rom[415][60] = 8'd38;
        rom[415][61] = -8'd4;
        rom[415][62] = 8'd19;
        rom[415][63] = -8'd3;
        rom[416][0] = -8'd24;
        rom[416][1] = 8'd41;
        rom[416][2] = 8'd9;
        rom[416][3] = -8'd11;
        rom[416][4] = 8'd3;
        rom[416][5] = 8'd23;
        rom[416][6] = 8'd22;
        rom[416][7] = 8'd17;
        rom[416][8] = -8'd17;
        rom[416][9] = -8'd5;
        rom[416][10] = -8'd4;
        rom[416][11] = 8'd50;
        rom[416][12] = -8'd21;
        rom[416][13] = -8'd62;
        rom[416][14] = -8'd35;
        rom[416][15] = -8'd32;
        rom[416][16] = -8'd27;
        rom[416][17] = -8'd13;
        rom[416][18] = -8'd39;
        rom[416][19] = -8'd41;
        rom[416][20] = -8'd1;
        rom[416][21] = 8'd13;
        rom[416][22] = 8'd1;
        rom[416][23] = -8'd9;
        rom[416][24] = 8'd15;
        rom[416][25] = -8'd2;
        rom[416][26] = -8'd6;
        rom[416][27] = 8'd1;
        rom[416][28] = 8'd13;
        rom[416][29] = 8'd47;
        rom[416][30] = -8'd19;
        rom[416][31] = 8'd20;
        rom[416][32] = -8'd41;
        rom[416][33] = -8'd23;
        rom[416][34] = 8'd0;
        rom[416][35] = 8'd7;
        rom[416][36] = -8'd14;
        rom[416][37] = -8'd7;
        rom[416][38] = -8'd18;
        rom[416][39] = 8'd26;
        rom[416][40] = -8'd50;
        rom[416][41] = 8'd14;
        rom[416][42] = 8'd11;
        rom[416][43] = 8'd11;
        rom[416][44] = -8'd9;
        rom[416][45] = -8'd6;
        rom[416][46] = -8'd34;
        rom[416][47] = 8'd24;
        rom[416][48] = 8'd66;
        rom[416][49] = -8'd15;
        rom[416][50] = 8'd7;
        rom[416][51] = 8'd1;
        rom[416][52] = -8'd36;
        rom[416][53] = -8'd45;
        rom[416][54] = 8'd35;
        rom[416][55] = -8'd37;
        rom[416][56] = -8'd6;
        rom[416][57] = -8'd57;
        rom[416][58] = 8'd13;
        rom[416][59] = -8'd45;
        rom[416][60] = 8'd14;
        rom[416][61] = 8'd9;
        rom[416][62] = 8'd28;
        rom[416][63] = 8'd12;
        rom[417][0] = 8'd29;
        rom[417][1] = -8'd18;
        rom[417][2] = -8'd30;
        rom[417][3] = 8'd11;
        rom[417][4] = 8'd27;
        rom[417][5] = 8'd4;
        rom[417][6] = -8'd15;
        rom[417][7] = 8'd18;
        rom[417][8] = -8'd19;
        rom[417][9] = -8'd6;
        rom[417][10] = 8'd10;
        rom[417][11] = 8'd20;
        rom[417][12] = -8'd21;
        rom[417][13] = -8'd4;
        rom[417][14] = -8'd39;
        rom[417][15] = 8'd34;
        rom[417][16] = 8'd22;
        rom[417][17] = -8'd32;
        rom[417][18] = 8'd1;
        rom[417][19] = 8'd23;
        rom[417][20] = -8'd5;
        rom[417][21] = -8'd36;
        rom[417][22] = -8'd18;
        rom[417][23] = -8'd5;
        rom[417][24] = 8'd48;
        rom[417][25] = -8'd8;
        rom[417][26] = 8'd6;
        rom[417][27] = 8'd11;
        rom[417][28] = 8'd34;
        rom[417][29] = -8'd36;
        rom[417][30] = -8'd20;
        rom[417][31] = 8'd19;
        rom[417][32] = 8'd32;
        rom[417][33] = -8'd19;
        rom[417][34] = -8'd41;
        rom[417][35] = -8'd52;
        rom[417][36] = -8'd9;
        rom[417][37] = -8'd2;
        rom[417][38] = -8'd96;
        rom[417][39] = 8'd19;
        rom[417][40] = -8'd21;
        rom[417][41] = 8'd0;
        rom[417][42] = 8'd37;
        rom[417][43] = 8'd9;
        rom[417][44] = -8'd24;
        rom[417][45] = -8'd20;
        rom[417][46] = 8'd19;
        rom[417][47] = 8'd28;
        rom[417][48] = -8'd50;
        rom[417][49] = -8'd16;
        rom[417][50] = 8'd18;
        rom[417][51] = -8'd13;
        rom[417][52] = -8'd2;
        rom[417][53] = -8'd50;
        rom[417][54] = -8'd25;
        rom[417][55] = -8'd31;
        rom[417][56] = 8'd35;
        rom[417][57] = 8'd20;
        rom[417][58] = -8'd8;
        rom[417][59] = 8'd17;
        rom[417][60] = 8'd66;
        rom[417][61] = -8'd1;
        rom[417][62] = 8'd24;
        rom[417][63] = 8'd30;
        rom[418][0] = -8'd14;
        rom[418][1] = 8'd10;
        rom[418][2] = 8'd12;
        rom[418][3] = 8'd4;
        rom[418][4] = -8'd5;
        rom[418][5] = -8'd8;
        rom[418][6] = -8'd30;
        rom[418][7] = 8'd45;
        rom[418][8] = -8'd6;
        rom[418][9] = 8'd26;
        rom[418][10] = 8'd34;
        rom[418][11] = 8'd7;
        rom[418][12] = -8'd39;
        rom[418][13] = 8'd22;
        rom[418][14] = 8'd5;
        rom[418][15] = -8'd12;
        rom[418][16] = -8'd17;
        rom[418][17] = 8'd10;
        rom[418][18] = 8'd17;
        rom[418][19] = -8'd3;
        rom[418][20] = -8'd5;
        rom[418][21] = 8'd0;
        rom[418][22] = 8'd6;
        rom[418][23] = 8'd48;
        rom[418][24] = 8'd5;
        rom[418][25] = 8'd0;
        rom[418][26] = 8'd47;
        rom[418][27] = -8'd68;
        rom[418][28] = -8'd5;
        rom[418][29] = -8'd2;
        rom[418][30] = -8'd10;
        rom[418][31] = -8'd20;
        rom[418][32] = -8'd32;
        rom[418][33] = -8'd3;
        rom[418][34] = -8'd19;
        rom[418][35] = -8'd20;
        rom[418][36] = 8'd16;
        rom[418][37] = 8'd5;
        rom[418][38] = 8'd4;
        rom[418][39] = 8'd15;
        rom[418][40] = 8'd5;
        rom[418][41] = -8'd23;
        rom[418][42] = -8'd14;
        rom[418][43] = -8'd27;
        rom[418][44] = 8'd25;
        rom[418][45] = 8'd22;
        rom[418][46] = -8'd14;
        rom[418][47] = -8'd10;
        rom[418][48] = 8'd45;
        rom[418][49] = -8'd40;
        rom[418][50] = -8'd11;
        rom[418][51] = 8'd48;
        rom[418][52] = 8'd20;
        rom[418][53] = 8'd17;
        rom[418][54] = -8'd11;
        rom[418][55] = 8'd20;
        rom[418][56] = 8'd18;
        rom[418][57] = 8'd23;
        rom[418][58] = -8'd38;
        rom[418][59] = 8'd2;
        rom[418][60] = -8'd16;
        rom[418][61] = 8'd27;
        rom[418][62] = -8'd13;
        rom[418][63] = 8'd21;
        rom[419][0] = -8'd23;
        rom[419][1] = -8'd50;
        rom[419][2] = -8'd50;
        rom[419][3] = -8'd13;
        rom[419][4] = -8'd17;
        rom[419][5] = -8'd30;
        rom[419][6] = 8'd26;
        rom[419][7] = -8'd19;
        rom[419][8] = -8'd3;
        rom[419][9] = 8'd10;
        rom[419][10] = -8'd49;
        rom[419][11] = -8'd7;
        rom[419][12] = -8'd44;
        rom[419][13] = -8'd4;
        rom[419][14] = -8'd20;
        rom[419][15] = -8'd15;
        rom[419][16] = -8'd7;
        rom[419][17] = -8'd4;
        rom[419][18] = -8'd57;
        rom[419][19] = -8'd9;
        rom[419][20] = -8'd1;
        rom[419][21] = -8'd32;
        rom[419][22] = -8'd44;
        rom[419][23] = -8'd12;
        rom[419][24] = -8'd9;
        rom[419][25] = 8'd6;
        rom[419][26] = -8'd23;
        rom[419][27] = 8'd34;
        rom[419][28] = -8'd17;
        rom[419][29] = -8'd14;
        rom[419][30] = -8'd38;
        rom[419][31] = 8'd14;
        rom[419][32] = 8'd14;
        rom[419][33] = -8'd30;
        rom[419][34] = -8'd1;
        rom[419][35] = -8'd13;
        rom[419][36] = 8'd15;
        rom[419][37] = -8'd79;
        rom[419][38] = -8'd19;
        rom[419][39] = 8'd9;
        rom[419][40] = -8'd29;
        rom[419][41] = 8'd16;
        rom[419][42] = -8'd34;
        rom[419][43] = 8'd0;
        rom[419][44] = -8'd15;
        rom[419][45] = -8'd14;
        rom[419][46] = -8'd40;
        rom[419][47] = -8'd9;
        rom[419][48] = -8'd21;
        rom[419][49] = 8'd12;
        rom[419][50] = -8'd52;
        rom[419][51] = 8'd5;
        rom[419][52] = -8'd39;
        rom[419][53] = 8'd8;
        rom[419][54] = 8'd17;
        rom[419][55] = -8'd34;
        rom[419][56] = -8'd2;
        rom[419][57] = -8'd65;
        rom[419][58] = -8'd27;
        rom[419][59] = -8'd30;
        rom[419][60] = -8'd14;
        rom[419][61] = -8'd3;
        rom[419][62] = -8'd17;
        rom[419][63] = 8'd3;
        rom[420][0] = -8'd5;
        rom[420][1] = 8'd13;
        rom[420][2] = 8'd7;
        rom[420][3] = -8'd36;
        rom[420][4] = -8'd34;
        rom[420][5] = 8'd43;
        rom[420][6] = 8'd25;
        rom[420][7] = -8'd84;
        rom[420][8] = -8'd26;
        rom[420][9] = -8'd18;
        rom[420][10] = 8'd46;
        rom[420][11] = 8'd12;
        rom[420][12] = -8'd12;
        rom[420][13] = -8'd5;
        rom[420][14] = -8'd21;
        rom[420][15] = -8'd26;
        rom[420][16] = -8'd27;
        rom[420][17] = -8'd13;
        rom[420][18] = 8'd13;
        rom[420][19] = 8'd4;
        rom[420][20] = -8'd12;
        rom[420][21] = -8'd9;
        rom[420][22] = 8'd12;
        rom[420][23] = -8'd47;
        rom[420][24] = -8'd53;
        rom[420][25] = -8'd24;
        rom[420][26] = 8'd14;
        rom[420][27] = -8'd40;
        rom[420][28] = 8'd29;
        rom[420][29] = 8'd6;
        rom[420][30] = 8'd6;
        rom[420][31] = -8'd50;
        rom[420][32] = 8'd0;
        rom[420][33] = 8'd14;
        rom[420][34] = 8'd2;
        rom[420][35] = -8'd4;
        rom[420][36] = -8'd14;
        rom[420][37] = -8'd17;
        rom[420][38] = -8'd9;
        rom[420][39] = -8'd10;
        rom[420][40] = 8'd8;
        rom[420][41] = 8'd13;
        rom[420][42] = 8'd31;
        rom[420][43] = -8'd22;
        rom[420][44] = 8'd2;
        rom[420][45] = -8'd49;
        rom[420][46] = -8'd17;
        rom[420][47] = 8'd44;
        rom[420][48] = -8'd24;
        rom[420][49] = 8'd14;
        rom[420][50] = 8'd5;
        rom[420][51] = -8'd6;
        rom[420][52] = -8'd22;
        rom[420][53] = 8'd11;
        rom[420][54] = -8'd15;
        rom[420][55] = -8'd13;
        rom[420][56] = 8'd16;
        rom[420][57] = -8'd37;
        rom[420][58] = 8'd25;
        rom[420][59] = -8'd23;
        rom[420][60] = -8'd37;
        rom[420][61] = 8'd8;
        rom[420][62] = 8'd24;
        rom[420][63] = 8'd44;
        rom[421][0] = -8'd16;
        rom[421][1] = 8'd8;
        rom[421][2] = -8'd52;
        rom[421][3] = 8'd29;
        rom[421][4] = -8'd43;
        rom[421][5] = -8'd15;
        rom[421][6] = 8'd40;
        rom[421][7] = -8'd79;
        rom[421][8] = 8'd34;
        rom[421][9] = 8'd57;
        rom[421][10] = -8'd72;
        rom[421][11] = 8'd8;
        rom[421][12] = -8'd44;
        rom[421][13] = -8'd5;
        rom[421][14] = -8'd30;
        rom[421][15] = 8'd9;
        rom[421][16] = 8'd24;
        rom[421][17] = -8'd54;
        rom[421][18] = -8'd18;
        rom[421][19] = -8'd51;
        rom[421][20] = 8'd8;
        rom[421][21] = 8'd3;
        rom[421][22] = -8'd40;
        rom[421][23] = -8'd3;
        rom[421][24] = -8'd4;
        rom[421][25] = 8'd57;
        rom[421][26] = 8'd27;
        rom[421][27] = 8'd12;
        rom[421][28] = 8'd27;
        rom[421][29] = 8'd18;
        rom[421][30] = 8'd14;
        rom[421][31] = 8'd24;
        rom[421][32] = 8'd9;
        rom[421][33] = 8'd17;
        rom[421][34] = -8'd1;
        rom[421][35] = -8'd1;
        rom[421][36] = -8'd45;
        rom[421][37] = 8'd9;
        rom[421][38] = -8'd35;
        rom[421][39] = -8'd22;
        rom[421][40] = 8'd2;
        rom[421][41] = 8'd28;
        rom[421][42] = -8'd41;
        rom[421][43] = -8'd72;
        rom[421][44] = 8'd34;
        rom[421][45] = -8'd26;
        rom[421][46] = -8'd35;
        rom[421][47] = 8'd3;
        rom[421][48] = 8'd4;
        rom[421][49] = 8'd17;
        rom[421][50] = 8'd23;
        rom[421][51] = 8'd7;
        rom[421][52] = 8'd21;
        rom[421][53] = -8'd30;
        rom[421][54] = -8'd8;
        rom[421][55] = -8'd21;
        rom[421][56] = -8'd10;
        rom[421][57] = -8'd45;
        rom[421][58] = 8'd17;
        rom[421][59] = -8'd61;
        rom[421][60] = 8'd9;
        rom[421][61] = -8'd37;
        rom[421][62] = 8'd35;
        rom[421][63] = 8'd46;
        rom[422][0] = -8'd13;
        rom[422][1] = -8'd12;
        rom[422][2] = 8'd3;
        rom[422][3] = 8'd21;
        rom[422][4] = 8'd25;
        rom[422][5] = -8'd26;
        rom[422][6] = -8'd97;
        rom[422][7] = -8'd7;
        rom[422][8] = -8'd40;
        rom[422][9] = -8'd5;
        rom[422][10] = 8'd6;
        rom[422][11] = 8'd23;
        rom[422][12] = 8'd36;
        rom[422][13] = 8'd17;
        rom[422][14] = 8'd10;
        rom[422][15] = -8'd5;
        rom[422][16] = 8'd26;
        rom[422][17] = -8'd58;
        rom[422][18] = -8'd69;
        rom[422][19] = -8'd35;
        rom[422][20] = -8'd14;
        rom[422][21] = -8'd16;
        rom[422][22] = 8'd6;
        rom[422][23] = 8'd32;
        rom[422][24] = 8'd5;
        rom[422][25] = -8'd41;
        rom[422][26] = -8'd19;
        rom[422][27] = -8'd5;
        rom[422][28] = -8'd19;
        rom[422][29] = 8'd24;
        rom[422][30] = 8'd5;
        rom[422][31] = -8'd16;
        rom[422][32] = 8'd19;
        rom[422][33] = -8'd13;
        rom[422][34] = 8'd13;
        rom[422][35] = -8'd37;
        rom[422][36] = -8'd16;
        rom[422][37] = 8'd6;
        rom[422][38] = 8'd38;
        rom[422][39] = 8'd1;
        rom[422][40] = 8'd16;
        rom[422][41] = 8'd35;
        rom[422][42] = 8'd17;
        rom[422][43] = 8'd11;
        rom[422][44] = -8'd17;
        rom[422][45] = 8'd0;
        rom[422][46] = 8'd22;
        rom[422][47] = -8'd13;
        rom[422][48] = -8'd45;
        rom[422][49] = -8'd16;
        rom[422][50] = 8'd14;
        rom[422][51] = -8'd32;
        rom[422][52] = -8'd4;
        rom[422][53] = -8'd6;
        rom[422][54] = -8'd28;
        rom[422][55] = -8'd33;
        rom[422][56] = 8'd5;
        rom[422][57] = 8'd25;
        rom[422][58] = 8'd37;
        rom[422][59] = 8'd36;
        rom[422][60] = -8'd29;
        rom[422][61] = -8'd10;
        rom[422][62] = 8'd2;
        rom[422][63] = 8'd14;
        rom[423][0] = -8'd31;
        rom[423][1] = -8'd4;
        rom[423][2] = -8'd31;
        rom[423][3] = 8'd4;
        rom[423][4] = 8'd2;
        rom[423][5] = -8'd11;
        rom[423][6] = -8'd2;
        rom[423][7] = -8'd3;
        rom[423][8] = 8'd2;
        rom[423][9] = -8'd6;
        rom[423][10] = -8'd17;
        rom[423][11] = 8'd8;
        rom[423][12] = -8'd4;
        rom[423][13] = -8'd15;
        rom[423][14] = -8'd6;
        rom[423][15] = -8'd33;
        rom[423][16] = -8'd39;
        rom[423][17] = 8'd30;
        rom[423][18] = 8'd12;
        rom[423][19] = 8'd0;
        rom[423][20] = 8'd3;
        rom[423][21] = -8'd10;
        rom[423][22] = 8'd0;
        rom[423][23] = -8'd61;
        rom[423][24] = 8'd2;
        rom[423][25] = 8'd10;
        rom[423][26] = 8'd32;
        rom[423][27] = 8'd23;
        rom[423][28] = 8'd2;
        rom[423][29] = 8'd12;
        rom[423][30] = 8'd23;
        rom[423][31] = 8'd0;
        rom[423][32] = -8'd18;
        rom[423][33] = 8'd1;
        rom[423][34] = 8'd16;
        rom[423][35] = 8'd10;
        rom[423][36] = 8'd13;
        rom[423][37] = 8'd2;
        rom[423][38] = -8'd12;
        rom[423][39] = 8'd26;
        rom[423][40] = -8'd2;
        rom[423][41] = -8'd2;
        rom[423][42] = -8'd6;
        rom[423][43] = -8'd9;
        rom[423][44] = -8'd12;
        rom[423][45] = -8'd12;
        rom[423][46] = -8'd12;
        rom[423][47] = -8'd39;
        rom[423][48] = -8'd22;
        rom[423][49] = 8'd6;
        rom[423][50] = 8'd16;
        rom[423][51] = -8'd25;
        rom[423][52] = -8'd4;
        rom[423][53] = -8'd24;
        rom[423][54] = 8'd26;
        rom[423][55] = 8'd9;
        rom[423][56] = 8'd20;
        rom[423][57] = 8'd63;
        rom[423][58] = -8'd30;
        rom[423][59] = 8'd14;
        rom[423][60] = -8'd38;
        rom[423][61] = 8'd8;
        rom[423][62] = 8'd30;
        rom[423][63] = -8'd32;
        rom[424][0] = 8'd9;
        rom[424][1] = 8'd22;
        rom[424][2] = 8'd14;
        rom[424][3] = 8'd5;
        rom[424][4] = 8'd12;
        rom[424][5] = 8'd2;
        rom[424][6] = 8'd12;
        rom[424][7] = -8'd2;
        rom[424][8] = 8'd32;
        rom[424][9] = 8'd40;
        rom[424][10] = -8'd108;
        rom[424][11] = -8'd5;
        rom[424][12] = 8'd7;
        rom[424][13] = 8'd15;
        rom[424][14] = 8'd13;
        rom[424][15] = -8'd31;
        rom[424][16] = -8'd31;
        rom[424][17] = 8'd25;
        rom[424][18] = 8'd25;
        rom[424][19] = 8'd7;
        rom[424][20] = -8'd4;
        rom[424][21] = -8'd23;
        rom[424][22] = 8'd1;
        rom[424][23] = -8'd10;
        rom[424][24] = 8'd27;
        rom[424][25] = -8'd14;
        rom[424][26] = -8'd21;
        rom[424][27] = -8'd4;
        rom[424][28] = 8'd23;
        rom[424][29] = 8'd6;
        rom[424][30] = -8'd17;
        rom[424][31] = -8'd20;
        rom[424][32] = 8'd17;
        rom[424][33] = -8'd14;
        rom[424][34] = -8'd19;
        rom[424][35] = 8'd23;
        rom[424][36] = 8'd2;
        rom[424][37] = 8'd2;
        rom[424][38] = 8'd34;
        rom[424][39] = -8'd9;
        rom[424][40] = 8'd16;
        rom[424][41] = -8'd22;
        rom[424][42] = 8'd10;
        rom[424][43] = 8'd26;
        rom[424][44] = 8'd23;
        rom[424][45] = 8'd28;
        rom[424][46] = -8'd5;
        rom[424][47] = -8'd28;
        rom[424][48] = 8'd40;
        rom[424][49] = -8'd24;
        rom[424][50] = 8'd10;
        rom[424][51] = -8'd15;
        rom[424][52] = -8'd27;
        rom[424][53] = 8'd40;
        rom[424][54] = 8'd9;
        rom[424][55] = -8'd17;
        rom[424][56] = 8'd13;
        rom[424][57] = -8'd5;
        rom[424][58] = -8'd5;
        rom[424][59] = -8'd30;
        rom[424][60] = 8'd20;
        rom[424][61] = -8'd22;
        rom[424][62] = 8'd38;
        rom[424][63] = 8'd12;
        rom[425][0] = -8'd66;
        rom[425][1] = 8'd54;
        rom[425][2] = -8'd22;
        rom[425][3] = 8'd6;
        rom[425][4] = -8'd22;
        rom[425][5] = -8'd50;
        rom[425][6] = 8'd36;
        rom[425][7] = -8'd66;
        rom[425][8] = 8'd11;
        rom[425][9] = 8'd9;
        rom[425][10] = -8'd76;
        rom[425][11] = -8'd56;
        rom[425][12] = -8'd9;
        rom[425][13] = -8'd3;
        rom[425][14] = 8'd0;
        rom[425][15] = -8'd20;
        rom[425][16] = -8'd7;
        rom[425][17] = -8'd38;
        rom[425][18] = -8'd20;
        rom[425][19] = -8'd13;
        rom[425][20] = 8'd6;
        rom[425][21] = -8'd26;
        rom[425][22] = -8'd12;
        rom[425][23] = -8'd82;
        rom[425][24] = 8'd12;
        rom[425][25] = 8'd14;
        rom[425][26] = 8'd18;
        rom[425][27] = 8'd9;
        rom[425][28] = -8'd7;
        rom[425][29] = 8'd14;
        rom[425][30] = -8'd36;
        rom[425][31] = 8'd17;
        rom[425][32] = -8'd8;
        rom[425][33] = -8'd22;
        rom[425][34] = 8'd28;
        rom[425][35] = -8'd50;
        rom[425][36] = 8'd61;
        rom[425][37] = -8'd16;
        rom[425][38] = -8'd35;
        rom[425][39] = -8'd35;
        rom[425][40] = 8'd8;
        rom[425][41] = 8'd20;
        rom[425][42] = -8'd29;
        rom[425][43] = 8'd1;
        rom[425][44] = 8'd19;
        rom[425][45] = -8'd93;
        rom[425][46] = -8'd16;
        rom[425][47] = -8'd91;
        rom[425][48] = -8'd38;
        rom[425][49] = 8'd15;
        rom[425][50] = 8'd28;
        rom[425][51] = 8'd23;
        rom[425][52] = 8'd23;
        rom[425][53] = -8'd39;
        rom[425][54] = -8'd41;
        rom[425][55] = 8'd5;
        rom[425][56] = -8'd26;
        rom[425][57] = 8'd37;
        rom[425][58] = -8'd19;
        rom[425][59] = 8'd4;
        rom[425][60] = 8'd13;
        rom[425][61] = 8'd23;
        rom[425][62] = -8'd24;
        rom[425][63] = -8'd7;
        rom[426][0] = 8'd14;
        rom[426][1] = 8'd1;
        rom[426][2] = -8'd28;
        rom[426][3] = 8'd36;
        rom[426][4] = 8'd5;
        rom[426][5] = 8'd4;
        rom[426][6] = 8'd3;
        rom[426][7] = -8'd3;
        rom[426][8] = -8'd15;
        rom[426][9] = 8'd3;
        rom[426][10] = -8'd9;
        rom[426][11] = 8'd22;
        rom[426][12] = 8'd7;
        rom[426][13] = -8'd24;
        rom[426][14] = -8'd3;
        rom[426][15] = 8'd6;
        rom[426][16] = -8'd47;
        rom[426][17] = -8'd41;
        rom[426][18] = 8'd11;
        rom[426][19] = 8'd12;
        rom[426][20] = -8'd2;
        rom[426][21] = 8'd36;
        rom[426][22] = 8'd11;
        rom[426][23] = 8'd4;
        rom[426][24] = 8'd2;
        rom[426][25] = -8'd109;
        rom[426][26] = 8'd14;
        rom[426][27] = 8'd53;
        rom[426][28] = 8'd19;
        rom[426][29] = -8'd20;
        rom[426][30] = -8'd12;
        rom[426][31] = 8'd11;
        rom[426][32] = 8'd25;
        rom[426][33] = 8'd31;
        rom[426][34] = -8'd7;
        rom[426][35] = -8'd13;
        rom[426][36] = -8'd28;
        rom[426][37] = -8'd5;
        rom[426][38] = 8'd5;
        rom[426][39] = 8'd12;
        rom[426][40] = 8'd6;
        rom[426][41] = 8'd28;
        rom[426][42] = 8'd12;
        rom[426][43] = -8'd33;
        rom[426][44] = -8'd33;
        rom[426][45] = 8'd7;
        rom[426][46] = 8'd13;
        rom[426][47] = -8'd20;
        rom[426][48] = 8'd19;
        rom[426][49] = -8'd16;
        rom[426][50] = 8'd1;
        rom[426][51] = -8'd36;
        rom[426][52] = -8'd41;
        rom[426][53] = 8'd11;
        rom[426][54] = -8'd19;
        rom[426][55] = -8'd13;
        rom[426][56] = -8'd32;
        rom[426][57] = 8'd42;
        rom[426][58] = -8'd4;
        rom[426][59] = 8'd23;
        rom[426][60] = 8'd13;
        rom[426][61] = 8'd46;
        rom[426][62] = -8'd34;
        rom[426][63] = -8'd22;
        rom[427][0] = 8'd16;
        rom[427][1] = -8'd6;
        rom[427][2] = 8'd5;
        rom[427][3] = -8'd46;
        rom[427][4] = -8'd7;
        rom[427][5] = 8'd12;
        rom[427][6] = -8'd3;
        rom[427][7] = -8'd11;
        rom[427][8] = -8'd24;
        rom[427][9] = 8'd20;
        rom[427][10] = -8'd7;
        rom[427][11] = 8'd49;
        rom[427][12] = 8'd24;
        rom[427][13] = -8'd39;
        rom[427][14] = 8'd18;
        rom[427][15] = -8'd3;
        rom[427][16] = 8'd28;
        rom[427][17] = -8'd25;
        rom[427][18] = 8'd6;
        rom[427][19] = 8'd14;
        rom[427][20] = -8'd9;
        rom[427][21] = 8'd26;
        rom[427][22] = -8'd6;
        rom[427][23] = 8'd7;
        rom[427][24] = -8'd17;
        rom[427][25] = 8'd13;
        rom[427][26] = 8'd19;
        rom[427][27] = 8'd44;
        rom[427][28] = 8'd7;
        rom[427][29] = -8'd3;
        rom[427][30] = 8'd24;
        rom[427][31] = 8'd35;
        rom[427][32] = -8'd7;
        rom[427][33] = 8'd9;
        rom[427][34] = 8'd10;
        rom[427][35] = -8'd4;
        rom[427][36] = 8'd20;
        rom[427][37] = -8'd46;
        rom[427][38] = 8'd25;
        rom[427][39] = -8'd26;
        rom[427][40] = -8'd15;
        rom[427][41] = 8'd26;
        rom[427][42] = 8'd17;
        rom[427][43] = -8'd12;
        rom[427][44] = 8'd27;
        rom[427][45] = 8'd1;
        rom[427][46] = -8'd19;
        rom[427][47] = -8'd28;
        rom[427][48] = 8'd0;
        rom[427][49] = 8'd2;
        rom[427][50] = 8'd41;
        rom[427][51] = -8'd7;
        rom[427][52] = -8'd21;
        rom[427][53] = -8'd10;
        rom[427][54] = -8'd19;
        rom[427][55] = 8'd46;
        rom[427][56] = -8'd2;
        rom[427][57] = -8'd9;
        rom[427][58] = 8'd14;
        rom[427][59] = -8'd8;
        rom[427][60] = -8'd11;
        rom[427][61] = -8'd20;
        rom[427][62] = 8'd23;
        rom[427][63] = 8'd15;
        rom[428][0] = -8'd23;
        rom[428][1] = 8'd2;
        rom[428][2] = -8'd68;
        rom[428][3] = 8'd45;
        rom[428][4] = 8'd21;
        rom[428][5] = -8'd20;
        rom[428][6] = -8'd16;
        rom[428][7] = 8'd1;
        rom[428][8] = -8'd25;
        rom[428][9] = 8'd17;
        rom[428][10] = 8'd19;
        rom[428][11] = 8'd3;
        rom[428][12] = 8'd6;
        rom[428][13] = -8'd13;
        rom[428][14] = -8'd13;
        rom[428][15] = -8'd20;
        rom[428][16] = 8'd1;
        rom[428][17] = 8'd7;
        rom[428][18] = -8'd17;
        rom[428][19] = -8'd39;
        rom[428][20] = -8'd12;
        rom[428][21] = 8'd29;
        rom[428][22] = 8'd4;
        rom[428][23] = -8'd22;
        rom[428][24] = -8'd13;
        rom[428][25] = 8'd0;
        rom[428][26] = 8'd8;
        rom[428][27] = -8'd13;
        rom[428][28] = 8'd5;
        rom[428][29] = -8'd83;
        rom[428][30] = 8'd20;
        rom[428][31] = -8'd29;
        rom[428][32] = -8'd28;
        rom[428][33] = -8'd8;
        rom[428][34] = 8'd22;
        rom[428][35] = -8'd26;
        rom[428][36] = -8'd41;
        rom[428][37] = -8'd8;
        rom[428][38] = -8'd22;
        rom[428][39] = 8'd12;
        rom[428][40] = 8'd46;
        rom[428][41] = -8'd43;
        rom[428][42] = -8'd2;
        rom[428][43] = -8'd32;
        rom[428][44] = -8'd10;
        rom[428][45] = -8'd3;
        rom[428][46] = -8'd34;
        rom[428][47] = 8'd5;
        rom[428][48] = -8'd42;
        rom[428][49] = 8'd19;
        rom[428][50] = -8'd23;
        rom[428][51] = 8'd40;
        rom[428][52] = 8'd24;
        rom[428][53] = 8'd17;
        rom[428][54] = -8'd1;
        rom[428][55] = 8'd31;
        rom[428][56] = 8'd1;
        rom[428][57] = 8'd14;
        rom[428][58] = 8'd4;
        rom[428][59] = 8'd4;
        rom[428][60] = 8'd13;
        rom[428][61] = -8'd11;
        rom[428][62] = 8'd9;
        rom[428][63] = 8'd16;
        rom[429][0] = 8'd1;
        rom[429][1] = 8'd10;
        rom[429][2] = -8'd30;
        rom[429][3] = -8'd5;
        rom[429][4] = 8'd22;
        rom[429][5] = -8'd81;
        rom[429][6] = -8'd25;
        rom[429][7] = -8'd83;
        rom[429][8] = 8'd34;
        rom[429][9] = 8'd13;
        rom[429][10] = -8'd19;
        rom[429][11] = 8'd40;
        rom[429][12] = 8'd3;
        rom[429][13] = 8'd3;
        rom[429][14] = -8'd8;
        rom[429][15] = -8'd16;
        rom[429][16] = 8'd5;
        rom[429][17] = -8'd20;
        rom[429][18] = -8'd28;
        rom[429][19] = -8'd26;
        rom[429][20] = 8'd2;
        rom[429][21] = 8'd7;
        rom[429][22] = -8'd32;
        rom[429][23] = -8'd54;
        rom[429][24] = -8'd43;
        rom[429][25] = -8'd21;
        rom[429][26] = -8'd40;
        rom[429][27] = -8'd45;
        rom[429][28] = -8'd32;
        rom[429][29] = -8'd11;
        rom[429][30] = -8'd1;
        rom[429][31] = -8'd61;
        rom[429][32] = 8'd26;
        rom[429][33] = 8'd27;
        rom[429][34] = 8'd60;
        rom[429][35] = 8'd5;
        rom[429][36] = -8'd60;
        rom[429][37] = 8'd19;
        rom[429][38] = -8'd9;
        rom[429][39] = 8'd5;
        rom[429][40] = -8'd36;
        rom[429][41] = 8'd21;
        rom[429][42] = -8'd43;
        rom[429][43] = -8'd21;
        rom[429][44] = -8'd21;
        rom[429][45] = -8'd51;
        rom[429][46] = -8'd60;
        rom[429][47] = 8'd71;
        rom[429][48] = 8'd20;
        rom[429][49] = 8'd11;
        rom[429][50] = -8'd16;
        rom[429][51] = -8'd28;
        rom[429][52] = -8'd23;
        rom[429][53] = -8'd3;
        rom[429][54] = 8'd20;
        rom[429][55] = -8'd3;
        rom[429][56] = 8'd9;
        rom[429][57] = -8'd18;
        rom[429][58] = -8'd8;
        rom[429][59] = -8'd16;
        rom[429][60] = 8'd31;
        rom[429][61] = 8'd1;
        rom[429][62] = -8'd9;
        rom[429][63] = 8'd37;
        rom[430][0] = -8'd16;
        rom[430][1] = -8'd38;
        rom[430][2] = 8'd1;
        rom[430][3] = 8'd17;
        rom[430][4] = 8'd7;
        rom[430][5] = 8'd3;
        rom[430][6] = 8'd17;
        rom[430][7] = 8'd3;
        rom[430][8] = 8'd28;
        rom[430][9] = -8'd3;
        rom[430][10] = -8'd18;
        rom[430][11] = 8'd32;
        rom[430][12] = -8'd44;
        rom[430][13] = -8'd47;
        rom[430][14] = -8'd7;
        rom[430][15] = -8'd30;
        rom[430][16] = -8'd128;
        rom[430][17] = -8'd33;
        rom[430][18] = -8'd22;
        rom[430][19] = 8'd17;
        rom[430][20] = 8'd1;
        rom[430][21] = 8'd13;
        rom[430][22] = -8'd22;
        rom[430][23] = -8'd43;
        rom[430][24] = 8'd3;
        rom[430][25] = 8'd41;
        rom[430][26] = 8'd20;
        rom[430][27] = -8'd40;
        rom[430][28] = 8'd12;
        rom[430][29] = -8'd12;
        rom[430][30] = -8'd9;
        rom[430][31] = -8'd40;
        rom[430][32] = 8'd26;
        rom[430][33] = -8'd34;
        rom[430][34] = -8'd14;
        rom[430][35] = 8'd23;
        rom[430][36] = 8'd40;
        rom[430][37] = -8'd109;
        rom[430][38] = -8'd10;
        rom[430][39] = 8'd7;
        rom[430][40] = -8'd22;
        rom[430][41] = -8'd14;
        rom[430][42] = -8'd15;
        rom[430][43] = 8'd1;
        rom[430][44] = -8'd49;
        rom[430][45] = -8'd48;
        rom[430][46] = -8'd15;
        rom[430][47] = -8'd41;
        rom[430][48] = -8'd21;
        rom[430][49] = 8'd16;
        rom[430][50] = -8'd48;
        rom[430][51] = 8'd5;
        rom[430][52] = -8'd10;
        rom[430][53] = 8'd17;
        rom[430][54] = -8'd6;
        rom[430][55] = 8'd18;
        rom[430][56] = -8'd9;
        rom[430][57] = 8'd28;
        rom[430][58] = -8'd2;
        rom[430][59] = -8'd77;
        rom[430][60] = 8'd14;
        rom[430][61] = 8'd14;
        rom[430][62] = 8'd28;
        rom[430][63] = 8'd6;
        rom[431][0] = -8'd23;
        rom[431][1] = 8'd52;
        rom[431][2] = -8'd61;
        rom[431][3] = -8'd1;
        rom[431][4] = 8'd10;
        rom[431][5] = 8'd6;
        rom[431][6] = 8'd2;
        rom[431][7] = 8'd68;
        rom[431][8] = -8'd47;
        rom[431][9] = 8'd8;
        rom[431][10] = 8'd0;
        rom[431][11] = 8'd11;
        rom[431][12] = 8'd1;
        rom[431][13] = -8'd6;
        rom[431][14] = 8'd25;
        rom[431][15] = -8'd28;
        rom[431][16] = -8'd13;
        rom[431][17] = 8'd17;
        rom[431][18] = -8'd12;
        rom[431][19] = 8'd22;
        rom[431][20] = 8'd8;
        rom[431][21] = 8'd35;
        rom[431][22] = 8'd46;
        rom[431][23] = 8'd41;
        rom[431][24] = 8'd30;
        rom[431][25] = -8'd5;
        rom[431][26] = -8'd2;
        rom[431][27] = 8'd8;
        rom[431][28] = 8'd44;
        rom[431][29] = -8'd33;
        rom[431][30] = -8'd7;
        rom[431][31] = 8'd5;
        rom[431][32] = 8'd40;
        rom[431][33] = 8'd14;
        rom[431][34] = 8'd37;
        rom[431][35] = 8'd11;
        rom[431][36] = -8'd4;
        rom[431][37] = 8'd51;
        rom[431][38] = -8'd15;
        rom[431][39] = 8'd17;
        rom[431][40] = -8'd39;
        rom[431][41] = -8'd11;
        rom[431][42] = 8'd42;
        rom[431][43] = 8'd8;
        rom[431][44] = 8'd11;
        rom[431][45] = -8'd9;
        rom[431][46] = -8'd33;
        rom[431][47] = 8'd12;
        rom[431][48] = 8'd30;
        rom[431][49] = 8'd15;
        rom[431][50] = -8'd49;
        rom[431][51] = 8'd28;
        rom[431][52] = 8'd5;
        rom[431][53] = 8'd41;
        rom[431][54] = -8'd22;
        rom[431][55] = -8'd33;
        rom[431][56] = 8'd13;
        rom[431][57] = 8'd57;
        rom[431][58] = 8'd1;
        rom[431][59] = -8'd42;
        rom[431][60] = 8'd10;
        rom[431][61] = -8'd27;
        rom[431][62] = 8'd1;
        rom[431][63] = 8'd33;
        rom[432][0] = 8'd40;
        rom[432][1] = 8'd4;
        rom[432][2] = -8'd45;
        rom[432][3] = 8'd22;
        rom[432][4] = -8'd22;
        rom[432][5] = 8'd8;
        rom[432][6] = 8'd15;
        rom[432][7] = 8'd1;
        rom[432][8] = 8'd20;
        rom[432][9] = -8'd11;
        rom[432][10] = 8'd11;
        rom[432][11] = -8'd4;
        rom[432][12] = -8'd19;
        rom[432][13] = -8'd30;
        rom[432][14] = -8'd37;
        rom[432][15] = 8'd3;
        rom[432][16] = 8'd28;
        rom[432][17] = 8'd17;
        rom[432][18] = 8'd15;
        rom[432][19] = 8'd29;
        rom[432][20] = -8'd7;
        rom[432][21] = 8'd22;
        rom[432][22] = -8'd19;
        rom[432][23] = 8'd49;
        rom[432][24] = 8'd24;
        rom[432][25] = -8'd2;
        rom[432][26] = 8'd2;
        rom[432][27] = 8'd12;
        rom[432][28] = 8'd44;
        rom[432][29] = -8'd5;
        rom[432][30] = -8'd6;
        rom[432][31] = 8'd46;
        rom[432][32] = 8'd32;
        rom[432][33] = 8'd54;
        rom[432][34] = -8'd33;
        rom[432][35] = -8'd22;
        rom[432][36] = 8'd27;
        rom[432][37] = -8'd63;
        rom[432][38] = 8'd10;
        rom[432][39] = 8'd1;
        rom[432][40] = -8'd11;
        rom[432][41] = -8'd44;
        rom[432][42] = -8'd1;
        rom[432][43] = 8'd21;
        rom[432][44] = 8'd29;
        rom[432][45] = -8'd2;
        rom[432][46] = 8'd2;
        rom[432][47] = 8'd28;
        rom[432][48] = 8'd6;
        rom[432][49] = -8'd4;
        rom[432][50] = -8'd43;
        rom[432][51] = -8'd17;
        rom[432][52] = -8'd33;
        rom[432][53] = -8'd1;
        rom[432][54] = -8'd22;
        rom[432][55] = 8'd6;
        rom[432][56] = -8'd9;
        rom[432][57] = -8'd2;
        rom[432][58] = 8'd38;
        rom[432][59] = 8'd7;
        rom[432][60] = -8'd42;
        rom[432][61] = 8'd5;
        rom[432][62] = -8'd2;
        rom[432][63] = -8'd5;
        rom[433][0] = -8'd27;
        rom[433][1] = 8'd28;
        rom[433][2] = -8'd11;
        rom[433][3] = 8'd4;
        rom[433][4] = -8'd3;
        rom[433][5] = -8'd35;
        rom[433][6] = -8'd5;
        rom[433][7] = 8'd14;
        rom[433][8] = 8'd10;
        rom[433][9] = 8'd1;
        rom[433][10] = 8'd14;
        rom[433][11] = 8'd38;
        rom[433][12] = 8'd36;
        rom[433][13] = 8'd37;
        rom[433][14] = 8'd14;
        rom[433][15] = -8'd13;
        rom[433][16] = -8'd72;
        rom[433][17] = -8'd29;
        rom[433][18] = -8'd19;
        rom[433][19] = 8'd13;
        rom[433][20] = 8'd3;
        rom[433][21] = -8'd43;
        rom[433][22] = 8'd30;
        rom[433][23] = -8'd3;
        rom[433][24] = 8'd5;
        rom[433][25] = -8'd7;
        rom[433][26] = -8'd21;
        rom[433][27] = -8'd43;
        rom[433][28] = 8'd8;
        rom[433][29] = 8'd21;
        rom[433][30] = 8'd12;
        rom[433][31] = -8'd18;
        rom[433][32] = 8'd29;
        rom[433][33] = -8'd4;
        rom[433][34] = -8'd17;
        rom[433][35] = 8'd46;
        rom[433][36] = 8'd36;
        rom[433][37] = -8'd22;
        rom[433][38] = 8'd7;
        rom[433][39] = -8'd65;
        rom[433][40] = 8'd6;
        rom[433][41] = 8'd12;
        rom[433][42] = 8'd9;
        rom[433][43] = -8'd24;
        rom[433][44] = 8'd18;
        rom[433][45] = 8'd10;
        rom[433][46] = 8'd50;
        rom[433][47] = 8'd17;
        rom[433][48] = -8'd32;
        rom[433][49] = 8'd44;
        rom[433][50] = 8'd12;
        rom[433][51] = -8'd24;
        rom[433][52] = -8'd22;
        rom[433][53] = 8'd14;
        rom[433][54] = -8'd36;
        rom[433][55] = -8'd36;
        rom[433][56] = 8'd27;
        rom[433][57] = 8'd47;
        rom[433][58] = -8'd11;
        rom[433][59] = -8'd17;
        rom[433][60] = 8'd38;
        rom[433][61] = 8'd32;
        rom[433][62] = 8'd10;
        rom[433][63] = 8'd22;
        rom[434][0] = 8'd4;
        rom[434][1] = -8'd6;
        rom[434][2] = 8'd29;
        rom[434][3] = 8'd11;
        rom[434][4] = 8'd20;
        rom[434][5] = -8'd5;
        rom[434][6] = -8'd19;
        rom[434][7] = 8'd19;
        rom[434][8] = -8'd27;
        rom[434][9] = 8'd26;
        rom[434][10] = -8'd36;
        rom[434][11] = 8'd1;
        rom[434][12] = -8'd15;
        rom[434][13] = 8'd19;
        rom[434][14] = -8'd58;
        rom[434][15] = 8'd8;
        rom[434][16] = -8'd45;
        rom[434][17] = -8'd17;
        rom[434][18] = 8'd26;
        rom[434][19] = -8'd25;
        rom[434][20] = -8'd9;
        rom[434][21] = -8'd20;
        rom[434][22] = 8'd10;
        rom[434][23] = -8'd33;
        rom[434][24] = -8'd11;
        rom[434][25] = -8'd16;
        rom[434][26] = 8'd3;
        rom[434][27] = 8'd70;
        rom[434][28] = 8'd9;
        rom[434][29] = 8'd18;
        rom[434][30] = 8'd4;
        rom[434][31] = -8'd59;
        rom[434][32] = 8'd4;
        rom[434][33] = -8'd38;
        rom[434][34] = 8'd41;
        rom[434][35] = 8'd16;
        rom[434][36] = -8'd1;
        rom[434][37] = -8'd53;
        rom[434][38] = -8'd53;
        rom[434][39] = -8'd36;
        rom[434][40] = 8'd15;
        rom[434][41] = 8'd8;
        rom[434][42] = -8'd8;
        rom[434][43] = 8'd12;
        rom[434][44] = 8'd29;
        rom[434][45] = -8'd60;
        rom[434][46] = 8'd4;
        rom[434][47] = 8'd2;
        rom[434][48] = -8'd15;
        rom[434][49] = -8'd17;
        rom[434][50] = 8'd15;
        rom[434][51] = -8'd33;
        rom[434][52] = 8'd10;
        rom[434][53] = -8'd21;
        rom[434][54] = -8'd27;
        rom[434][55] = -8'd8;
        rom[434][56] = -8'd18;
        rom[434][57] = -8'd41;
        rom[434][58] = -8'd38;
        rom[434][59] = -8'd27;
        rom[434][60] = 8'd10;
        rom[434][61] = -8'd56;
        rom[434][62] = -8'd31;
        rom[434][63] = 8'd7;
        rom[435][0] = 8'd25;
        rom[435][1] = -8'd27;
        rom[435][2] = 8'd15;
        rom[435][3] = 8'd27;
        rom[435][4] = -8'd43;
        rom[435][5] = -8'd4;
        rom[435][6] = -8'd4;
        rom[435][7] = 8'd7;
        rom[435][8] = -8'd7;
        rom[435][9] = 8'd15;
        rom[435][10] = 8'd8;
        rom[435][11] = -8'd25;
        rom[435][12] = 8'd24;
        rom[435][13] = -8'd11;
        rom[435][14] = -8'd31;
        rom[435][15] = -8'd11;
        rom[435][16] = -8'd22;
        rom[435][17] = 8'd3;
        rom[435][18] = 8'd2;
        rom[435][19] = -8'd1;
        rom[435][20] = 8'd2;
        rom[435][21] = -8'd8;
        rom[435][22] = -8'd17;
        rom[435][23] = -8'd16;
        rom[435][24] = 8'd3;
        rom[435][25] = -8'd37;
        rom[435][26] = -8'd1;
        rom[435][27] = 8'd2;
        rom[435][28] = 8'd23;
        rom[435][29] = -8'd9;
        rom[435][30] = -8'd70;
        rom[435][31] = 8'd15;
        rom[435][32] = -8'd42;
        rom[435][33] = -8'd31;
        rom[435][34] = 8'd3;
        rom[435][35] = -8'd29;
        rom[435][36] = -8'd21;
        rom[435][37] = -8'd25;
        rom[435][38] = -8'd1;
        rom[435][39] = -8'd21;
        rom[435][40] = -8'd23;
        rom[435][41] = -8'd4;
        rom[435][42] = -8'd64;
        rom[435][43] = -8'd28;
        rom[435][44] = 8'd6;
        rom[435][45] = 8'd8;
        rom[435][46] = -8'd6;
        rom[435][47] = 8'd9;
        rom[435][48] = 8'd2;
        rom[435][49] = -8'd7;
        rom[435][50] = 8'd1;
        rom[435][51] = 8'd18;
        rom[435][52] = -8'd6;
        rom[435][53] = -8'd31;
        rom[435][54] = 8'd30;
        rom[435][55] = -8'd20;
        rom[435][56] = -8'd18;
        rom[435][57] = 8'd22;
        rom[435][58] = 8'd45;
        rom[435][59] = 8'd10;
        rom[435][60] = -8'd26;
        rom[435][61] = 8'd6;
        rom[435][62] = 8'd27;
        rom[435][63] = 8'd43;
        rom[436][0] = 8'd33;
        rom[436][1] = -8'd2;
        rom[436][2] = -8'd26;
        rom[436][3] = -8'd9;
        rom[436][4] = 8'd27;
        rom[436][5] = 8'd16;
        rom[436][6] = -8'd103;
        rom[436][7] = 8'd14;
        rom[436][8] = -8'd12;
        rom[436][9] = -8'd15;
        rom[436][10] = 8'd49;
        rom[436][11] = 8'd32;
        rom[436][12] = -8'd38;
        rom[436][13] = 8'd12;
        rom[436][14] = -8'd12;
        rom[436][15] = -8'd1;
        rom[436][16] = -8'd21;
        rom[436][17] = 8'd39;
        rom[436][18] = 8'd9;
        rom[436][19] = -8'd42;
        rom[436][20] = -8'd13;
        rom[436][21] = 8'd24;
        rom[436][22] = -8'd43;
        rom[436][23] = -8'd2;
        rom[436][24] = -8'd43;
        rom[436][25] = 8'd1;
        rom[436][26] = -8'd2;
        rom[436][27] = 8'd38;
        rom[436][28] = 8'd36;
        rom[436][29] = -8'd28;
        rom[436][30] = -8'd5;
        rom[436][31] = -8'd12;
        rom[436][32] = 8'd22;
        rom[436][33] = 8'd80;
        rom[436][34] = 8'd13;
        rom[436][35] = 8'd13;
        rom[436][36] = -8'd13;
        rom[436][37] = 8'd53;
        rom[436][38] = 8'd18;
        rom[436][39] = 8'd40;
        rom[436][40] = 8'd18;
        rom[436][41] = -8'd17;
        rom[436][42] = -8'd26;
        rom[436][43] = 8'd9;
        rom[436][44] = 8'd6;
        rom[436][45] = 8'd23;
        rom[436][46] = 8'd31;
        rom[436][47] = -8'd2;
        rom[436][48] = 8'd15;
        rom[436][49] = 8'd15;
        rom[436][50] = 8'd19;
        rom[436][51] = -8'd28;
        rom[436][52] = 8'd26;
        rom[436][53] = 8'd8;
        rom[436][54] = 8'd4;
        rom[436][55] = -8'd33;
        rom[436][56] = 8'd41;
        rom[436][57] = -8'd33;
        rom[436][58] = 8'd38;
        rom[436][59] = -8'd34;
        rom[436][60] = -8'd53;
        rom[436][61] = -8'd15;
        rom[436][62] = 8'd29;
        rom[436][63] = -8'd29;
        rom[437][0] = 8'd31;
        rom[437][1] = 8'd18;
        rom[437][2] = 8'd8;
        rom[437][3] = 8'd15;
        rom[437][4] = 8'd16;
        rom[437][5] = 8'd2;
        rom[437][6] = -8'd19;
        rom[437][7] = 8'd28;
        rom[437][8] = 8'd9;
        rom[437][9] = -8'd42;
        rom[437][10] = -8'd28;
        rom[437][11] = -8'd39;
        rom[437][12] = -8'd14;
        rom[437][13] = -8'd4;
        rom[437][14] = -8'd17;
        rom[437][15] = -8'd1;
        rom[437][16] = -8'd13;
        rom[437][17] = -8'd6;
        rom[437][18] = 8'd3;
        rom[437][19] = -8'd4;
        rom[437][20] = -8'd3;
        rom[437][21] = -8'd16;
        rom[437][22] = -8'd34;
        rom[437][23] = 8'd13;
        rom[437][24] = -8'd38;
        rom[437][25] = 8'd13;
        rom[437][26] = -8'd28;
        rom[437][27] = -8'd49;
        rom[437][28] = -8'd16;
        rom[437][29] = 8'd25;
        rom[437][30] = 8'd23;
        rom[437][31] = -8'd43;
        rom[437][32] = -8'd3;
        rom[437][33] = 8'd10;
        rom[437][34] = -8'd2;
        rom[437][35] = -8'd9;
        rom[437][36] = 8'd1;
        rom[437][37] = -8'd17;
        rom[437][38] = -8'd40;
        rom[437][39] = -8'd44;
        rom[437][40] = 8'd10;
        rom[437][41] = -8'd20;
        rom[437][42] = -8'd28;
        rom[437][43] = 8'd26;
        rom[437][44] = -8'd5;
        rom[437][45] = -8'd23;
        rom[437][46] = -8'd24;
        rom[437][47] = 8'd13;
        rom[437][48] = 8'd1;
        rom[437][49] = -8'd34;
        rom[437][50] = -8'd36;
        rom[437][51] = -8'd43;
        rom[437][52] = 8'd9;
        rom[437][53] = 8'd29;
        rom[437][54] = -8'd4;
        rom[437][55] = -8'd28;
        rom[437][56] = -8'd39;
        rom[437][57] = -8'd14;
        rom[437][58] = -8'd16;
        rom[437][59] = 8'd50;
        rom[437][60] = -8'd24;
        rom[437][61] = 8'd0;
        rom[437][62] = -8'd7;
        rom[437][63] = -8'd28;
        rom[438][0] = -8'd1;
        rom[438][1] = 8'd4;
        rom[438][2] = 8'd4;
        rom[438][3] = 8'd4;
        rom[438][4] = 8'd2;
        rom[438][5] = -8'd6;
        rom[438][6] = -8'd7;
        rom[438][7] = -8'd13;
        rom[438][8] = 8'd11;
        rom[438][9] = -8'd5;
        rom[438][10] = 8'd2;
        rom[438][11] = 8'd5;
        rom[438][12] = -8'd3;
        rom[438][13] = -8'd3;
        rom[438][14] = -8'd4;
        rom[438][15] = -8'd8;
        rom[438][16] = 8'd14;
        rom[438][17] = -8'd1;
        rom[438][18] = -8'd8;
        rom[438][19] = 8'd9;
        rom[438][20] = 8'd3;
        rom[438][21] = 8'd0;
        rom[438][22] = -8'd5;
        rom[438][23] = 8'd7;
        rom[438][24] = -8'd9;
        rom[438][25] = -8'd10;
        rom[438][26] = -8'd2;
        rom[438][27] = 8'd7;
        rom[438][28] = 8'd9;
        rom[438][29] = 8'd1;
        rom[438][30] = 8'd5;
        rom[438][31] = -8'd6;
        rom[438][32] = -8'd1;
        rom[438][33] = 8'd5;
        rom[438][34] = -8'd8;
        rom[438][35] = 8'd5;
        rom[438][36] = -8'd2;
        rom[438][37] = -8'd7;
        rom[438][38] = -8'd4;
        rom[438][39] = -8'd4;
        rom[438][40] = 8'd5;
        rom[438][41] = -8'd3;
        rom[438][42] = 8'd9;
        rom[438][43] = -8'd8;
        rom[438][44] = -8'd4;
        rom[438][45] = -8'd2;
        rom[438][46] = 8'd6;
        rom[438][47] = 8'd14;
        rom[438][48] = -8'd2;
        rom[438][49] = 8'd3;
        rom[438][50] = 8'd4;
        rom[438][51] = -8'd2;
        rom[438][52] = 8'd7;
        rom[438][53] = 8'd10;
        rom[438][54] = -8'd4;
        rom[438][55] = 8'd5;
        rom[438][56] = 8'd0;
        rom[438][57] = -8'd5;
        rom[438][58] = 8'd2;
        rom[438][59] = 8'd0;
        rom[438][60] = 8'd9;
        rom[438][61] = 8'd4;
        rom[438][62] = 8'd12;
        rom[438][63] = 8'd5;
        rom[439][0] = -8'd14;
        rom[439][1] = 8'd10;
        rom[439][2] = -8'd22;
        rom[439][3] = 8'd2;
        rom[439][4] = -8'd1;
        rom[439][5] = 8'd3;
        rom[439][6] = -8'd85;
        rom[439][7] = 8'd6;
        rom[439][8] = -8'd33;
        rom[439][9] = 8'd21;
        rom[439][10] = 8'd11;
        rom[439][11] = -8'd19;
        rom[439][12] = 8'd9;
        rom[439][13] = 8'd2;
        rom[439][14] = -8'd39;
        rom[439][15] = -8'd16;
        rom[439][16] = 8'd12;
        rom[439][17] = -8'd18;
        rom[439][18] = -8'd25;
        rom[439][19] = -8'd38;
        rom[439][20] = 8'd2;
        rom[439][21] = 8'd9;
        rom[439][22] = -8'd34;
        rom[439][23] = -8'd20;
        rom[439][24] = -8'd15;
        rom[439][25] = 8'd22;
        rom[439][26] = 8'd26;
        rom[439][27] = -8'd48;
        rom[439][28] = 8'd10;
        rom[439][29] = -8'd34;
        rom[439][30] = 8'd12;
        rom[439][31] = -8'd17;
        rom[439][32] = -8'd54;
        rom[439][33] = 8'd17;
        rom[439][34] = 8'd26;
        rom[439][35] = -8'd35;
        rom[439][36] = -8'd1;
        rom[439][37] = 8'd7;
        rom[439][38] = -8'd5;
        rom[439][39] = 8'd21;
        rom[439][40] = 8'd35;
        rom[439][41] = -8'd31;
        rom[439][42] = -8'd26;
        rom[439][43] = -8'd37;
        rom[439][44] = 8'd18;
        rom[439][45] = -8'd4;
        rom[439][46] = -8'd3;
        rom[439][47] = -8'd25;
        rom[439][48] = -8'd24;
        rom[439][49] = -8'd12;
        rom[439][50] = -8'd13;
        rom[439][51] = -8'd3;
        rom[439][52] = -8'd22;
        rom[439][53] = -8'd3;
        rom[439][54] = -8'd31;
        rom[439][55] = -8'd42;
        rom[439][56] = 8'd16;
        rom[439][57] = 8'd25;
        rom[439][58] = 8'd8;
        rom[439][59] = 8'd14;
        rom[439][60] = -8'd91;
        rom[439][61] = 8'd0;
        rom[439][62] = 8'd1;
        rom[439][63] = 8'd27;
        rom[440][0] = -8'd5;
        rom[440][1] = -8'd6;
        rom[440][2] = 8'd14;
        rom[440][3] = 8'd38;
        rom[440][4] = -8'd47;
        rom[440][5] = -8'd25;
        rom[440][6] = -8'd18;
        rom[440][7] = -8'd1;
        rom[440][8] = 8'd7;
        rom[440][9] = -8'd24;
        rom[440][10] = 8'd22;
        rom[440][11] = 8'd20;
        rom[440][12] = 8'd19;
        rom[440][13] = -8'd2;
        rom[440][14] = 8'd28;
        rom[440][15] = -8'd6;
        rom[440][16] = 8'd6;
        rom[440][17] = 8'd11;
        rom[440][18] = -8'd40;
        rom[440][19] = 8'd16;
        rom[440][20] = -8'd6;
        rom[440][21] = 8'd39;
        rom[440][22] = 8'd8;
        rom[440][23] = 8'd56;
        rom[440][24] = 8'd47;
        rom[440][25] = -8'd30;
        rom[440][26] = -8'd4;
        rom[440][27] = -8'd23;
        rom[440][28] = 8'd34;
        rom[440][29] = -8'd19;
        rom[440][30] = -8'd4;
        rom[440][31] = -8'd80;
        rom[440][32] = 8'd26;
        rom[440][33] = -8'd18;
        rom[440][34] = -8'd14;
        rom[440][35] = -8'd21;
        rom[440][36] = -8'd8;
        rom[440][37] = -8'd26;
        rom[440][38] = -8'd7;
        rom[440][39] = 8'd5;
        rom[440][40] = 8'd24;
        rom[440][41] = -8'd1;
        rom[440][42] = -8'd4;
        rom[440][43] = -8'd27;
        rom[440][44] = 8'd0;
        rom[440][45] = 8'd7;
        rom[440][46] = -8'd52;
        rom[440][47] = 8'd5;
        rom[440][48] = 8'd31;
        rom[440][49] = 8'd10;
        rom[440][50] = -8'd27;
        rom[440][51] = -8'd17;
        rom[440][52] = -8'd2;
        rom[440][53] = 8'd0;
        rom[440][54] = 8'd21;
        rom[440][55] = 8'd10;
        rom[440][56] = -8'd4;
        rom[440][57] = 8'd11;
        rom[440][58] = 8'd9;
        rom[440][59] = -8'd3;
        rom[440][60] = 8'd4;
        rom[440][61] = 8'd4;
        rom[440][62] = 8'd19;
        rom[440][63] = 8'd36;
        rom[441][0] = 8'd9;
        rom[441][1] = 8'd33;
        rom[441][2] = -8'd2;
        rom[441][3] = 8'd18;
        rom[441][4] = -8'd5;
        rom[441][5] = 8'd8;
        rom[441][6] = -8'd23;
        rom[441][7] = 8'd1;
        rom[441][8] = -8'd25;
        rom[441][9] = 8'd1;
        rom[441][10] = 8'd14;
        rom[441][11] = -8'd22;
        rom[441][12] = 8'd33;
        rom[441][13] = -8'd6;
        rom[441][14] = -8'd5;
        rom[441][15] = 8'd3;
        rom[441][16] = -8'd4;
        rom[441][17] = 8'd16;
        rom[441][18] = -8'd8;
        rom[441][19] = -8'd12;
        rom[441][20] = -8'd7;
        rom[441][21] = -8'd25;
        rom[441][22] = -8'd69;
        rom[441][23] = 8'd47;
        rom[441][24] = -8'd8;
        rom[441][25] = -8'd15;
        rom[441][26] = -8'd5;
        rom[441][27] = 8'd38;
        rom[441][28] = 8'd13;
        rom[441][29] = -8'd16;
        rom[441][30] = -8'd40;
        rom[441][31] = -8'd12;
        rom[441][32] = -8'd15;
        rom[441][33] = -8'd10;
        rom[441][34] = 8'd50;
        rom[441][35] = 8'd2;
        rom[441][36] = 8'd19;
        rom[441][37] = 8'd24;
        rom[441][38] = -8'd10;
        rom[441][39] = -8'd32;
        rom[441][40] = -8'd27;
        rom[441][41] = -8'd58;
        rom[441][42] = 8'd0;
        rom[441][43] = -8'd34;
        rom[441][44] = -8'd10;
        rom[441][45] = -8'd64;
        rom[441][46] = 8'd37;
        rom[441][47] = -8'd48;
        rom[441][48] = -8'd75;
        rom[441][49] = -8'd13;
        rom[441][50] = 8'd23;
        rom[441][51] = -8'd14;
        rom[441][52] = 8'd28;
        rom[441][53] = -8'd74;
        rom[441][54] = -8'd38;
        rom[441][55] = 8'd28;
        rom[441][56] = -8'd7;
        rom[441][57] = -8'd7;
        rom[441][58] = 8'd37;
        rom[441][59] = 8'd17;
        rom[441][60] = 8'd11;
        rom[441][61] = 8'd28;
        rom[441][62] = 8'd35;
        rom[441][63] = -8'd14;
        rom[442][0] = 8'd26;
        rom[442][1] = 8'd23;
        rom[442][2] = -8'd11;
        rom[442][3] = -8'd1;
        rom[442][4] = -8'd24;
        rom[442][5] = -8'd34;
        rom[442][6] = -8'd20;
        rom[442][7] = -8'd80;
        rom[442][8] = 8'd21;
        rom[442][9] = -8'd27;
        rom[442][10] = 8'd64;
        rom[442][11] = -8'd18;
        rom[442][12] = -8'd25;
        rom[442][13] = 8'd6;
        rom[442][14] = 8'd12;
        rom[442][15] = 8'd27;
        rom[442][16] = 8'd34;
        rom[442][17] = 8'd12;
        rom[442][18] = -8'd17;
        rom[442][19] = 8'd42;
        rom[442][20] = 8'd2;
        rom[442][21] = -8'd38;
        rom[442][22] = -8'd25;
        rom[442][23] = -8'd6;
        rom[442][24] = 8'd4;
        rom[442][25] = 8'd0;
        rom[442][26] = 8'd9;
        rom[442][27] = -8'd36;
        rom[442][28] = 8'd18;
        rom[442][29] = -8'd11;
        rom[442][30] = -8'd28;
        rom[442][31] = 8'd18;
        rom[442][32] = 8'd21;
        rom[442][33] = 8'd10;
        rom[442][34] = 8'd26;
        rom[442][35] = 8'd0;
        rom[442][36] = -8'd1;
        rom[442][37] = 8'd7;
        rom[442][38] = -8'd64;
        rom[442][39] = -8'd30;
        rom[442][40] = -8'd12;
        rom[442][41] = 8'd7;
        rom[442][42] = -8'd5;
        rom[442][43] = 8'd23;
        rom[442][44] = -8'd10;
        rom[442][45] = 8'd15;
        rom[442][46] = 8'd44;
        rom[442][47] = 8'd35;
        rom[442][48] = -8'd31;
        rom[442][49] = 8'd16;
        rom[442][50] = -8'd46;
        rom[442][51] = -8'd2;
        rom[442][52] = 8'd59;
        rom[442][53] = 8'd10;
        rom[442][54] = -8'd17;
        rom[442][55] = 8'd38;
        rom[442][56] = 8'd19;
        rom[442][57] = 8'd43;
        rom[442][58] = -8'd45;
        rom[442][59] = -8'd17;
        rom[442][60] = 8'd16;
        rom[442][61] = -8'd18;
        rom[442][62] = -8'd62;
        rom[442][63] = -8'd11;
        rom[443][0] = 8'd7;
        rom[443][1] = -8'd25;
        rom[443][2] = -8'd34;
        rom[443][3] = -8'd50;
        rom[443][4] = 8'd1;
        rom[443][5] = 8'd4;
        rom[443][6] = -8'd5;
        rom[443][7] = -8'd12;
        rom[443][8] = -8'd33;
        rom[443][9] = 8'd7;
        rom[443][10] = -8'd1;
        rom[443][11] = 8'd14;
        rom[443][12] = -8'd3;
        rom[443][13] = 8'd13;
        rom[443][14] = -8'd3;
        rom[443][15] = -8'd35;
        rom[443][16] = 8'd24;
        rom[443][17] = -8'd59;
        rom[443][18] = -8'd25;
        rom[443][19] = -8'd32;
        rom[443][20] = 8'd3;
        rom[443][21] = -8'd63;
        rom[443][22] = 8'd39;
        rom[443][23] = 8'd32;
        rom[443][24] = -8'd1;
        rom[443][25] = -8'd2;
        rom[443][26] = -8'd4;
        rom[443][27] = -8'd53;
        rom[443][28] = 8'd6;
        rom[443][29] = 8'd14;
        rom[443][30] = -8'd2;
        rom[443][31] = -8'd5;
        rom[443][32] = -8'd40;
        rom[443][33] = 8'd12;
        rom[443][34] = -8'd1;
        rom[443][35] = 8'd29;
        rom[443][36] = -8'd59;
        rom[443][37] = -8'd2;
        rom[443][38] = -8'd4;
        rom[443][39] = 8'd0;
        rom[443][40] = 8'd6;
        rom[443][41] = -8'd38;
        rom[443][42] = 8'd3;
        rom[443][43] = 8'd2;
        rom[443][44] = -8'd16;
        rom[443][45] = -8'd14;
        rom[443][46] = -8'd31;
        rom[443][47] = 8'd30;
        rom[443][48] = -8'd8;
        rom[443][49] = 8'd40;
        rom[443][50] = -8'd21;
        rom[443][51] = 8'd31;
        rom[443][52] = -8'd9;
        rom[443][53] = 8'd0;
        rom[443][54] = -8'd24;
        rom[443][55] = -8'd73;
        rom[443][56] = 8'd24;
        rom[443][57] = -8'd9;
        rom[443][58] = -8'd22;
        rom[443][59] = -8'd14;
        rom[443][60] = 8'd4;
        rom[443][61] = -8'd57;
        rom[443][62] = 8'd2;
        rom[443][63] = 8'd17;
        rom[444][0] = 8'd21;
        rom[444][1] = -8'd2;
        rom[444][2] = 8'd5;
        rom[444][3] = -8'd6;
        rom[444][4] = 8'd6;
        rom[444][5] = -8'd47;
        rom[444][6] = 8'd4;
        rom[444][7] = -8'd15;
        rom[444][8] = 8'd2;
        rom[444][9] = -8'd37;
        rom[444][10] = -8'd41;
        rom[444][11] = 8'd14;
        rom[444][12] = -8'd30;
        rom[444][13] = -8'd40;
        rom[444][14] = -8'd36;
        rom[444][15] = 8'd10;
        rom[444][16] = 8'd31;
        rom[444][17] = 8'd7;
        rom[444][18] = -8'd19;
        rom[444][19] = 8'd16;
        rom[444][20] = 8'd0;
        rom[444][21] = 8'd18;
        rom[444][22] = -8'd17;
        rom[444][23] = -8'd34;
        rom[444][24] = 8'd37;
        rom[444][25] = -8'd8;
        rom[444][26] = -8'd25;
        rom[444][27] = -8'd23;
        rom[444][28] = 8'd16;
        rom[444][29] = -8'd5;
        rom[444][30] = -8'd13;
        rom[444][31] = -8'd3;
        rom[444][32] = 8'd1;
        rom[444][33] = 8'd14;
        rom[444][34] = 8'd2;
        rom[444][35] = -8'd1;
        rom[444][36] = 8'd23;
        rom[444][37] = -8'd38;
        rom[444][38] = -8'd20;
        rom[444][39] = 8'd21;
        rom[444][40] = 8'd25;
        rom[444][41] = 8'd16;
        rom[444][42] = 8'd7;
        rom[444][43] = 8'd21;
        rom[444][44] = 8'd12;
        rom[444][45] = -8'd29;
        rom[444][46] = 8'd25;
        rom[444][47] = 8'd31;
        rom[444][48] = 8'd15;
        rom[444][49] = -8'd29;
        rom[444][50] = 8'd39;
        rom[444][51] = 8'd14;
        rom[444][52] = 8'd1;
        rom[444][53] = -8'd58;
        rom[444][54] = 8'd36;
        rom[444][55] = -8'd27;
        rom[444][56] = 8'd0;
        rom[444][57] = -8'd3;
        rom[444][58] = -8'd5;
        rom[444][59] = -8'd46;
        rom[444][60] = -8'd3;
        rom[444][61] = -8'd5;
        rom[444][62] = 8'd46;
        rom[444][63] = 8'd17;
        rom[445][0] = -8'd35;
        rom[445][1] = 8'd9;
        rom[445][2] = -8'd3;
        rom[445][3] = 8'd7;
        rom[445][4] = -8'd2;
        rom[445][5] = -8'd2;
        rom[445][6] = -8'd76;
        rom[445][7] = -8'd5;
        rom[445][8] = -8'd41;
        rom[445][9] = -8'd27;
        rom[445][10] = 8'd10;
        rom[445][11] = -8'd20;
        rom[445][12] = 8'd51;
        rom[445][13] = 8'd17;
        rom[445][14] = 8'd34;
        rom[445][15] = -8'd9;
        rom[445][16] = -8'd52;
        rom[445][17] = -8'd70;
        rom[445][18] = -8'd17;
        rom[445][19] = 8'd28;
        rom[445][20] = -8'd3;
        rom[445][21] = -8'd15;
        rom[445][22] = 8'd12;
        rom[445][23] = 8'd16;
        rom[445][24] = -8'd14;
        rom[445][25] = -8'd51;
        rom[445][26] = 8'd33;
        rom[445][27] = -8'd2;
        rom[445][28] = -8'd10;
        rom[445][29] = -8'd27;
        rom[445][30] = 8'd1;
        rom[445][31] = -8'd41;
        rom[445][32] = 8'd16;
        rom[445][33] = -8'd40;
        rom[445][34] = 8'd16;
        rom[445][35] = 8'd6;
        rom[445][36] = -8'd11;
        rom[445][37] = -8'd43;
        rom[445][38] = 8'd16;
        rom[445][39] = -8'd4;
        rom[445][40] = 8'd7;
        rom[445][41] = -8'd4;
        rom[445][42] = 8'd9;
        rom[445][43] = 8'd14;
        rom[445][44] = 8'd31;
        rom[445][45] = -8'd39;
        rom[445][46] = -8'd1;
        rom[445][47] = -8'd15;
        rom[445][48] = 8'd13;
        rom[445][49] = 8'd42;
        rom[445][50] = 8'd19;
        rom[445][51] = 8'd6;
        rom[445][52] = 8'd0;
        rom[445][53] = -8'd3;
        rom[445][54] = -8'd25;
        rom[445][55] = 8'd9;
        rom[445][56] = 8'd22;
        rom[445][57] = 8'd2;
        rom[445][58] = -8'd27;
        rom[445][59] = 8'd10;
        rom[445][60] = 8'd15;
        rom[445][61] = -8'd5;
        rom[445][62] = -8'd5;
        rom[445][63] = 8'd11;
        rom[446][0] = 8'd17;
        rom[446][1] = -8'd1;
        rom[446][2] = 8'd5;
        rom[446][3] = 8'd7;
        rom[446][4] = -8'd44;
        rom[446][5] = 8'd21;
        rom[446][6] = -8'd5;
        rom[446][7] = -8'd3;
        rom[446][8] = -8'd24;
        rom[446][9] = 8'd2;
        rom[446][10] = 8'd20;
        rom[446][11] = 8'd53;
        rom[446][12] = -8'd37;
        rom[446][13] = 8'd20;
        rom[446][14] = -8'd50;
        rom[446][15] = 8'd55;
        rom[446][16] = 8'd1;
        rom[446][17] = -8'd12;
        rom[446][18] = -8'd8;
        rom[446][19] = -8'd22;
        rom[446][20] = 8'd5;
        rom[446][21] = 8'd31;
        rom[446][22] = 8'd29;
        rom[446][23] = 8'd12;
        rom[446][24] = 8'd21;
        rom[446][25] = -8'd5;
        rom[446][26] = -8'd16;
        rom[446][27] = -8'd5;
        rom[446][28] = -8'd49;
        rom[446][29] = 8'd9;
        rom[446][30] = -8'd81;
        rom[446][31] = 8'd15;
        rom[446][32] = 8'd15;
        rom[446][33] = 8'd28;
        rom[446][34] = -8'd7;
        rom[446][35] = -8'd47;
        rom[446][36] = -8'd32;
        rom[446][37] = -8'd61;
        rom[446][38] = -8'd36;
        rom[446][39] = 8'd20;
        rom[446][40] = 8'd19;
        rom[446][41] = -8'd19;
        rom[446][42] = 8'd30;
        rom[446][43] = 8'd22;
        rom[446][44] = 8'd13;
        rom[446][45] = -8'd16;
        rom[446][46] = 8'd32;
        rom[446][47] = 8'd23;
        rom[446][48] = -8'd59;
        rom[446][49] = -8'd63;
        rom[446][50] = 8'd40;
        rom[446][51] = 8'd43;
        rom[446][52] = 8'd1;
        rom[446][53] = -8'd44;
        rom[446][54] = -8'd13;
        rom[446][55] = -8'd25;
        rom[446][56] = -8'd23;
        rom[446][57] = 8'd12;
        rom[446][58] = 8'd9;
        rom[446][59] = 8'd1;
        rom[446][60] = 8'd23;
        rom[446][61] = -8'd65;
        rom[446][62] = 8'd10;
        rom[446][63] = 8'd25;
        rom[447][0] = -8'd12;
        rom[447][1] = -8'd3;
        rom[447][2] = -8'd3;
        rom[447][3] = 8'd1;
        rom[447][4] = 8'd13;
        rom[447][5] = 8'd1;
        rom[447][6] = 8'd3;
        rom[447][7] = -8'd2;
        rom[447][8] = 8'd22;
        rom[447][9] = 8'd9;
        rom[447][10] = -8'd18;
        rom[447][11] = 8'd24;
        rom[447][12] = -8'd57;
        rom[447][13] = 8'd4;
        rom[447][14] = -8'd13;
        rom[447][15] = 8'd18;
        rom[447][16] = -8'd34;
        rom[447][17] = -8'd13;
        rom[447][18] = -8'd1;
        rom[447][19] = -8'd7;
        rom[447][20] = 8'd0;
        rom[447][21] = -8'd33;
        rom[447][22] = 8'd46;
        rom[447][23] = -8'd12;
        rom[447][24] = 8'd20;
        rom[447][25] = -8'd49;
        rom[447][26] = 8'd13;
        rom[447][27] = -8'd23;
        rom[447][28] = -8'd20;
        rom[447][29] = -8'd24;
        rom[447][30] = -8'd82;
        rom[447][31] = -8'd25;
        rom[447][32] = -8'd15;
        rom[447][33] = -8'd1;
        rom[447][34] = -8'd23;
        rom[447][35] = 8'd23;
        rom[447][36] = 8'd11;
        rom[447][37] = 8'd55;
        rom[447][38] = -8'd35;
        rom[447][39] = 8'd23;
        rom[447][40] = -8'd24;
        rom[447][41] = 8'd33;
        rom[447][42] = -8'd6;
        rom[447][43] = 8'd1;
        rom[447][44] = 8'd15;
        rom[447][45] = -8'd39;
        rom[447][46] = -8'd25;
        rom[447][47] = -8'd63;
        rom[447][48] = -8'd8;
        rom[447][49] = -8'd4;
        rom[447][50] = -8'd9;
        rom[447][51] = -8'd4;
        rom[447][52] = 8'd10;
        rom[447][53] = 8'd29;
        rom[447][54] = -8'd36;
        rom[447][55] = 8'd29;
        rom[447][56] = -8'd29;
        rom[447][57] = -8'd10;
        rom[447][58] = -8'd23;
        rom[447][59] = -8'd26;
        rom[447][60] = 8'd2;
        rom[447][61] = -8'd10;
        rom[447][62] = 8'd16;
        rom[447][63] = -8'd56;
        rom[448][0] = 8'd5;
        rom[448][1] = -8'd6;
        rom[448][2] = -8'd21;
        rom[448][3] = -8'd3;
        rom[448][4] = -8'd26;
        rom[448][5] = 8'd12;
        rom[448][6] = -8'd6;
        rom[448][7] = 8'd24;
        rom[448][8] = -8'd31;
        rom[448][9] = 8'd24;
        rom[448][10] = -8'd7;
        rom[448][11] = 8'd24;
        rom[448][12] = -8'd22;
        rom[448][13] = -8'd8;
        rom[448][14] = -8'd23;
        rom[448][15] = 8'd17;
        rom[448][16] = 8'd9;
        rom[448][17] = 8'd50;
        rom[448][18] = -8'd4;
        rom[448][19] = 8'd24;
        rom[448][20] = 8'd3;
        rom[448][21] = -8'd2;
        rom[448][22] = -8'd89;
        rom[448][23] = 8'd16;
        rom[448][24] = 8'd6;
        rom[448][25] = 8'd1;
        rom[448][26] = -8'd20;
        rom[448][27] = -8'd27;
        rom[448][28] = 8'd41;
        rom[448][29] = -8'd3;
        rom[448][30] = 8'd29;
        rom[448][31] = -8'd7;
        rom[448][32] = -8'd23;
        rom[448][33] = 8'd18;
        rom[448][34] = 8'd14;
        rom[448][35] = -8'd45;
        rom[448][36] = -8'd36;
        rom[448][37] = -8'd24;
        rom[448][38] = -8'd18;
        rom[448][39] = 8'd20;
        rom[448][40] = -8'd36;
        rom[448][41] = 8'd3;
        rom[448][42] = -8'd5;
        rom[448][43] = -8'd36;
        rom[448][44] = -8'd24;
        rom[448][45] = 8'd20;
        rom[448][46] = 8'd4;
        rom[448][47] = -8'd65;
        rom[448][48] = 8'd1;
        rom[448][49] = -8'd18;
        rom[448][50] = -8'd21;
        rom[448][51] = -8'd64;
        rom[448][52] = 8'd12;
        rom[448][53] = -8'd2;
        rom[448][54] = -8'd4;
        rom[448][55] = -8'd1;
        rom[448][56] = 8'd10;
        rom[448][57] = -8'd7;
        rom[448][58] = -8'd32;
        rom[448][59] = 8'd19;
        rom[448][60] = -8'd17;
        rom[448][61] = -8'd57;
        rom[448][62] = -8'd35;
        rom[448][63] = 8'd23;
        rom[449][0] = -8'd33;
        rom[449][1] = -8'd67;
        rom[449][2] = -8'd24;
        rom[449][3] = -8'd7;
        rom[449][4] = -8'd61;
        rom[449][5] = -8'd23;
        rom[449][6] = -8'd53;
        rom[449][7] = -8'd24;
        rom[449][8] = -8'd21;
        rom[449][9] = -8'd40;
        rom[449][10] = -8'd47;
        rom[449][11] = -8'd7;
        rom[449][12] = -8'd42;
        rom[449][13] = -8'd12;
        rom[449][14] = -8'd26;
        rom[449][15] = 8'd2;
        rom[449][16] = -8'd13;
        rom[449][17] = -8'd84;
        rom[449][18] = -8'd24;
        rom[449][19] = -8'd51;
        rom[449][20] = -8'd4;
        rom[449][21] = -8'd20;
        rom[449][22] = -8'd50;
        rom[449][23] = -8'd25;
        rom[449][24] = -8'd11;
        rom[449][25] = -8'd9;
        rom[449][26] = -8'd5;
        rom[449][27] = -8'd29;
        rom[449][28] = 8'd30;
        rom[449][29] = -8'd17;
        rom[449][30] = -8'd20;
        rom[449][31] = -8'd5;
        rom[449][32] = -8'd9;
        rom[449][33] = 8'd26;
        rom[449][34] = -8'd3;
        rom[449][35] = 8'd5;
        rom[449][36] = -8'd16;
        rom[449][37] = -8'd17;
        rom[449][38] = 8'd1;
        rom[449][39] = 8'd16;
        rom[449][40] = 8'd50;
        rom[449][41] = -8'd22;
        rom[449][42] = 8'd6;
        rom[449][43] = -8'd30;
        rom[449][44] = 8'd20;
        rom[449][45] = -8'd9;
        rom[449][46] = -8'd33;
        rom[449][47] = 8'd59;
        rom[449][48] = -8'd8;
        rom[449][49] = 8'd13;
        rom[449][50] = -8'd10;
        rom[449][51] = -8'd12;
        rom[449][52] = -8'd76;
        rom[449][53] = -8'd1;
        rom[449][54] = -8'd56;
        rom[449][55] = 8'd5;
        rom[449][56] = 8'd9;
        rom[449][57] = 8'd11;
        rom[449][58] = -8'd8;
        rom[449][59] = -8'd23;
        rom[449][60] = -8'd36;
        rom[449][61] = -8'd3;
        rom[449][62] = -8'd1;
        rom[449][63] = 8'd8;
        rom[450][0] = -8'd20;
        rom[450][1] = 8'd3;
        rom[450][2] = -8'd52;
        rom[450][3] = -8'd50;
        rom[450][4] = -8'd77;
        rom[450][5] = -8'd6;
        rom[450][6] = -8'd34;
        rom[450][7] = 8'd18;
        rom[450][8] = -8'd68;
        rom[450][9] = 8'd14;
        rom[450][10] = 8'd2;
        rom[450][11] = -8'd29;
        rom[450][12] = 8'd19;
        rom[450][13] = -8'd64;
        rom[450][14] = -8'd14;
        rom[450][15] = -8'd6;
        rom[450][16] = 8'd4;
        rom[450][17] = -8'd4;
        rom[450][18] = 8'd30;
        rom[450][19] = -8'd18;
        rom[450][20] = -8'd1;
        rom[450][21] = 8'd13;
        rom[450][22] = -8'd104;
        rom[450][23] = -8'd18;
        rom[450][24] = -8'd46;
        rom[450][25] = 8'd2;
        rom[450][26] = 8'd9;
        rom[450][27] = 8'd7;
        rom[450][28] = 8'd21;
        rom[450][29] = 8'd7;
        rom[450][30] = 8'd14;
        rom[450][31] = -8'd46;
        rom[450][32] = 8'd15;
        rom[450][33] = -8'd14;
        rom[450][34] = -8'd17;
        rom[450][35] = -8'd33;
        rom[450][36] = 8'd16;
        rom[450][37] = -8'd16;
        rom[450][38] = 8'd8;
        rom[450][39] = -8'd11;
        rom[450][40] = -8'd13;
        rom[450][41] = -8'd31;
        rom[450][42] = -8'd67;
        rom[450][43] = 8'd25;
        rom[450][44] = 8'd7;
        rom[450][45] = -8'd16;
        rom[450][46] = -8'd39;
        rom[450][47] = 8'd19;
        rom[450][48] = -8'd70;
        rom[450][49] = -8'd8;
        rom[450][50] = -8'd20;
        rom[450][51] = -8'd17;
        rom[450][52] = 8'd9;
        rom[450][53] = -8'd50;
        rom[450][54] = -8'd52;
        rom[450][55] = 8'd12;
        rom[450][56] = -8'd13;
        rom[450][57] = -8'd22;
        rom[450][58] = 8'd4;
        rom[450][59] = -8'd1;
        rom[450][60] = 8'd1;
        rom[450][61] = 8'd12;
        rom[450][62] = 8'd21;
        rom[450][63] = -8'd37;
        rom[451][0] = 8'd27;
        rom[451][1] = 8'd37;
        rom[451][2] = -8'd38;
        rom[451][3] = 8'd11;
        rom[451][4] = 8'd11;
        rom[451][5] = 8'd33;
        rom[451][6] = -8'd3;
        rom[451][7] = 8'd50;
        rom[451][8] = -8'd6;
        rom[451][9] = 8'd29;
        rom[451][10] = -8'd23;
        rom[451][11] = -8'd14;
        rom[451][12] = -8'd42;
        rom[451][13] = -8'd21;
        rom[451][14] = 8'd44;
        rom[451][15] = 8'd21;
        rom[451][16] = -8'd52;
        rom[451][17] = 8'd36;
        rom[451][18] = 8'd3;
        rom[451][19] = -8'd3;
        rom[451][20] = -8'd3;
        rom[451][21] = -8'd16;
        rom[451][22] = -8'd2;
        rom[451][23] = 8'd9;
        rom[451][24] = 8'd1;
        rom[451][25] = -8'd25;
        rom[451][26] = 8'd36;
        rom[451][27] = -8'd23;
        rom[451][28] = 8'd17;
        rom[451][29] = 8'd3;
        rom[451][30] = 8'd6;
        rom[451][31] = 8'd26;
        rom[451][32] = -8'd24;
        rom[451][33] = 8'd19;
        rom[451][34] = 8'd11;
        rom[451][35] = -8'd28;
        rom[451][36] = -8'd6;
        rom[451][37] = -8'd16;
        rom[451][38] = -8'd61;
        rom[451][39] = 8'd32;
        rom[451][40] = 8'd6;
        rom[451][41] = 8'd5;
        rom[451][42] = -8'd5;
        rom[451][43] = -8'd27;
        rom[451][44] = -8'd24;
        rom[451][45] = -8'd16;
        rom[451][46] = -8'd63;
        rom[451][47] = -8'd50;
        rom[451][48] = 8'd24;
        rom[451][49] = -8'd8;
        rom[451][50] = -8'd25;
        rom[451][51] = -8'd3;
        rom[451][52] = 8'd21;
        rom[451][53] = 8'd15;
        rom[451][54] = -8'd13;
        rom[451][55] = -8'd43;
        rom[451][56] = 8'd9;
        rom[451][57] = -8'd79;
        rom[451][58] = 8'd30;
        rom[451][59] = 8'd12;
        rom[451][60] = 8'd2;
        rom[451][61] = -8'd25;
        rom[451][62] = -8'd28;
        rom[451][63] = 8'd3;
        rom[452][0] = -8'd25;
        rom[452][1] = -8'd27;
        rom[452][2] = -8'd71;
        rom[452][3] = 8'd1;
        rom[452][4] = -8'd24;
        rom[452][5] = -8'd27;
        rom[452][6] = -8'd10;
        rom[452][7] = -8'd5;
        rom[452][8] = 8'd0;
        rom[452][9] = -8'd19;
        rom[452][10] = -8'd22;
        rom[452][11] = 8'd18;
        rom[452][12] = -8'd7;
        rom[452][13] = -8'd2;
        rom[452][14] = -8'd10;
        rom[452][15] = -8'd21;
        rom[452][16] = 8'd31;
        rom[452][17] = -8'd8;
        rom[452][18] = 8'd4;
        rom[452][19] = 8'd15;
        rom[452][20] = 8'd7;
        rom[452][21] = -8'd41;
        rom[452][22] = -8'd12;
        rom[452][23] = -8'd28;
        rom[452][24] = -8'd21;
        rom[452][25] = -8'd6;
        rom[452][26] = -8'd29;
        rom[452][27] = 8'd0;
        rom[452][28] = -8'd17;
        rom[452][29] = -8'd9;
        rom[452][30] = -8'd46;
        rom[452][31] = -8'd40;
        rom[452][32] = 8'd32;
        rom[452][33] = -8'd11;
        rom[452][34] = 8'd8;
        rom[452][35] = 8'd4;
        rom[452][36] = 8'd0;
        rom[452][37] = -8'd22;
        rom[452][38] = -8'd8;
        rom[452][39] = -8'd43;
        rom[452][40] = -8'd6;
        rom[452][41] = 8'd16;
        rom[452][42] = -8'd32;
        rom[452][43] = -8'd57;
        rom[452][44] = -8'd5;
        rom[452][45] = -8'd5;
        rom[452][46] = -8'd25;
        rom[452][47] = -8'd52;
        rom[452][48] = -8'd7;
        rom[452][49] = -8'd39;
        rom[452][50] = -8'd34;
        rom[452][51] = -8'd12;
        rom[452][52] = -8'd77;
        rom[452][53] = -8'd15;
        rom[452][54] = -8'd6;
        rom[452][55] = -8'd10;
        rom[452][56] = -8'd31;
        rom[452][57] = -8'd12;
        rom[452][58] = -8'd2;
        rom[452][59] = -8'd35;
        rom[452][60] = 8'd48;
        rom[452][61] = 8'd11;
        rom[452][62] = 8'd4;
        rom[452][63] = -8'd14;
        rom[453][0] = 8'd6;
        rom[453][1] = 8'd5;
        rom[453][2] = -8'd6;
        rom[453][3] = 8'd4;
        rom[453][4] = -8'd8;
        rom[453][5] = 8'd7;
        rom[453][6] = 8'd8;
        rom[453][7] = 8'd4;
        rom[453][8] = 8'd1;
        rom[453][9] = 8'd2;
        rom[453][10] = 8'd5;
        rom[453][11] = 8'd0;
        rom[453][12] = -8'd8;
        rom[453][13] = 8'd7;
        rom[453][14] = -8'd5;
        rom[453][15] = 8'd2;
        rom[453][16] = 8'd4;
        rom[453][17] = -8'd2;
        rom[453][18] = -8'd3;
        rom[453][19] = 8'd7;
        rom[453][20] = -8'd5;
        rom[453][21] = 8'd1;
        rom[453][22] = -8'd15;
        rom[453][23] = 8'd8;
        rom[453][24] = 8'd7;
        rom[453][25] = 8'd7;
        rom[453][26] = 8'd12;
        rom[453][27] = -8'd4;
        rom[453][28] = -8'd1;
        rom[453][29] = 8'd12;
        rom[453][30] = 8'd1;
        rom[453][31] = -8'd3;
        rom[453][32] = 8'd5;
        rom[453][33] = 8'd1;
        rom[453][34] = -8'd3;
        rom[453][35] = 8'd2;
        rom[453][36] = -8'd8;
        rom[453][37] = 8'd1;
        rom[453][38] = -8'd5;
        rom[453][39] = -8'd1;
        rom[453][40] = 8'd11;
        rom[453][41] = -8'd13;
        rom[453][42] = 8'd10;
        rom[453][43] = -8'd3;
        rom[453][44] = 8'd6;
        rom[453][45] = 8'd0;
        rom[453][46] = 8'd2;
        rom[453][47] = -8'd2;
        rom[453][48] = -8'd5;
        rom[453][49] = 8'd1;
        rom[453][50] = 8'd0;
        rom[453][51] = 8'd1;
        rom[453][52] = -8'd6;
        rom[453][53] = -8'd7;
        rom[453][54] = 8'd6;
        rom[453][55] = 8'd3;
        rom[453][56] = 8'd5;
        rom[453][57] = -8'd12;
        rom[453][58] = 8'd16;
        rom[453][59] = 8'd8;
        rom[453][60] = 8'd3;
        rom[453][61] = 8'd0;
        rom[453][62] = 8'd4;
        rom[453][63] = 8'd1;
        rom[454][0] = 8'd28;
        rom[454][1] = -8'd16;
        rom[454][2] = 8'd21;
        rom[454][3] = -8'd17;
        rom[454][4] = -8'd90;
        rom[454][5] = 8'd33;
        rom[454][6] = -8'd17;
        rom[454][7] = 8'd0;
        rom[454][8] = 8'd6;
        rom[454][9] = 8'd23;
        rom[454][10] = 8'd7;
        rom[454][11] = 8'd51;
        rom[454][12] = -8'd33;
        rom[454][13] = 8'd12;
        rom[454][14] = -8'd37;
        rom[454][15] = -8'd1;
        rom[454][16] = -8'd50;
        rom[454][17] = 8'd43;
        rom[454][18] = 8'd32;
        rom[454][19] = -8'd52;
        rom[454][20] = -8'd5;
        rom[454][21] = 8'd5;
        rom[454][22] = 8'd3;
        rom[454][23] = 8'd57;
        rom[454][24] = -8'd8;
        rom[454][25] = 8'd11;
        rom[454][26] = 8'd33;
        rom[454][27] = -8'd51;
        rom[454][28] = 8'd15;
        rom[454][29] = 8'd24;
        rom[454][30] = 8'd22;
        rom[454][31] = 8'd17;
        rom[454][32] = -8'd26;
        rom[454][33] = -8'd10;
        rom[454][34] = 8'd34;
        rom[454][35] = 8'd0;
        rom[454][36] = -8'd29;
        rom[454][37] = -8'd3;
        rom[454][38] = 8'd23;
        rom[454][39] = -8'd10;
        rom[454][40] = 8'd15;
        rom[454][41] = -8'd30;
        rom[454][42] = 8'd28;
        rom[454][43] = -8'd16;
        rom[454][44] = -8'd6;
        rom[454][45] = 8'd14;
        rom[454][46] = 8'd1;
        rom[454][47] = 8'd6;
        rom[454][48] = 8'd31;
        rom[454][49] = -8'd19;
        rom[454][50] = -8'd2;
        rom[454][51] = -8'd2;
        rom[454][52] = -8'd18;
        rom[454][53] = -8'd50;
        rom[454][54] = 8'd44;
        rom[454][55] = -8'd9;
        rom[454][56] = 8'd33;
        rom[454][57] = 8'd23;
        rom[454][58] = 8'd26;
        rom[454][59] = -8'd23;
        rom[454][60] = -8'd24;
        rom[454][61] = -8'd35;
        rom[454][62] = 8'd21;
        rom[454][63] = 8'd4;
        rom[455][0] = 8'd27;
        rom[455][1] = -8'd24;
        rom[455][2] = -8'd21;
        rom[455][3] = 8'd0;
        rom[455][4] = -8'd10;
        rom[455][5] = 8'd26;
        rom[455][6] = 8'd6;
        rom[455][7] = 8'd1;
        rom[455][8] = 8'd8;
        rom[455][9] = -8'd17;
        rom[455][10] = -8'd2;
        rom[455][11] = -8'd47;
        rom[455][12] = -8'd61;
        rom[455][13] = 8'd37;
        rom[455][14] = -8'd13;
        rom[455][15] = 8'd29;
        rom[455][16] = -8'd10;
        rom[455][17] = -8'd22;
        rom[455][18] = -8'd28;
        rom[455][19] = 8'd15;
        rom[455][20] = 8'd6;
        rom[455][21] = 8'd29;
        rom[455][22] = 8'd23;
        rom[455][23] = 8'd16;
        rom[455][24] = -8'd1;
        rom[455][25] = 8'd4;
        rom[455][26] = -8'd3;
        rom[455][27] = 8'd2;
        rom[455][28] = 8'd41;
        rom[455][29] = -8'd8;
        rom[455][30] = -8'd79;
        rom[455][31] = -8'd80;
        rom[455][32] = 8'd32;
        rom[455][33] = 8'd5;
        rom[455][34] = 8'd19;
        rom[455][35] = -8'd1;
        rom[455][36] = 8'd6;
        rom[455][37] = -8'd3;
        rom[455][38] = -8'd2;
        rom[455][39] = 8'd0;
        rom[455][40] = 8'd8;
        rom[455][41] = -8'd8;
        rom[455][42] = 8'd23;
        rom[455][43] = 8'd27;
        rom[455][44] = -8'd15;
        rom[455][45] = -8'd1;
        rom[455][46] = 8'd45;
        rom[455][47] = -8'd7;
        rom[455][48] = -8'd11;
        rom[455][49] = -8'd9;
        rom[455][50] = -8'd16;
        rom[455][51] = 8'd15;
        rom[455][52] = -8'd34;
        rom[455][53] = 8'd5;
        rom[455][54] = -8'd56;
        rom[455][55] = -8'd3;
        rom[455][56] = 8'd0;
        rom[455][57] = -8'd12;
        rom[455][58] = -8'd21;
        rom[455][59] = -8'd16;
        rom[455][60] = 8'd5;
        rom[455][61] = -8'd11;
        rom[455][62] = 8'd15;
        rom[455][63] = 8'd5;
        rom[456][0] = -8'd3;
        rom[456][1] = 8'd10;
        rom[456][2] = 8'd4;
        rom[456][3] = -8'd10;
        rom[456][4] = 8'd17;
        rom[456][5] = -8'd26;
        rom[456][6] = -8'd18;
        rom[456][7] = -8'd50;
        rom[456][8] = -8'd1;
        rom[456][9] = -8'd31;
        rom[456][10] = 8'd14;
        rom[456][11] = -8'd25;
        rom[456][12] = -8'd25;
        rom[456][13] = -8'd27;
        rom[456][14] = -8'd4;
        rom[456][15] = -8'd20;
        rom[456][16] = -8'd36;
        rom[456][17] = 8'd5;
        rom[456][18] = -8'd12;
        rom[456][19] = -8'd19;
        rom[456][20] = -8'd6;
        rom[456][21] = -8'd27;
        rom[456][22] = -8'd18;
        rom[456][23] = 8'd15;
        rom[456][24] = -8'd18;
        rom[456][25] = -8'd23;
        rom[456][26] = -8'd30;
        rom[456][27] = -8'd14;
        rom[456][28] = 8'd6;
        rom[456][29] = 8'd0;
        rom[456][30] = -8'd64;
        rom[456][31] = 8'd10;
        rom[456][32] = -8'd6;
        rom[456][33] = 8'd9;
        rom[456][34] = -8'd1;
        rom[456][35] = 8'd4;
        rom[456][36] = -8'd4;
        rom[456][37] = -8'd16;
        rom[456][38] = -8'd15;
        rom[456][39] = 8'd18;
        rom[456][40] = -8'd49;
        rom[456][41] = -8'd8;
        rom[456][42] = -8'd11;
        rom[456][43] = 8'd33;
        rom[456][44] = -8'd12;
        rom[456][45] = -8'd10;
        rom[456][46] = -8'd6;
        rom[456][47] = -8'd37;
        rom[456][48] = -8'd37;
        rom[456][49] = 8'd13;
        rom[456][50] = -8'd30;
        rom[456][51] = -8'd24;
        rom[456][52] = -8'd8;
        rom[456][53] = -8'd34;
        rom[456][54] = -8'd18;
        rom[456][55] = 8'd21;
        rom[456][56] = 8'd1;
        rom[456][57] = -8'd12;
        rom[456][58] = 8'd3;
        rom[456][59] = -8'd22;
        rom[456][60] = 8'd11;
        rom[456][61] = -8'd37;
        rom[456][62] = -8'd12;
        rom[456][63] = -8'd36;
        rom[457][0] = -8'd28;
        rom[457][1] = -8'd37;
        rom[457][2] = 8'd17;
        rom[457][3] = -8'd2;
        rom[457][4] = -8'd2;
        rom[457][5] = 8'd10;
        rom[457][6] = 8'd11;
        rom[457][7] = 8'd4;
        rom[457][8] = 8'd16;
        rom[457][9] = -8'd59;
        rom[457][10] = -8'd38;
        rom[457][11] = -8'd15;
        rom[457][12] = 8'd32;
        rom[457][13] = 8'd2;
        rom[457][14] = -8'd3;
        rom[457][15] = -8'd11;
        rom[457][16] = -8'd46;
        rom[457][17] = -8'd27;
        rom[457][18] = -8'd4;
        rom[457][19] = -8'd12;
        rom[457][20] = -8'd5;
        rom[457][21] = 8'd24;
        rom[457][22] = 8'd58;
        rom[457][23] = 8'd0;
        rom[457][24] = 8'd1;
        rom[457][25] = -8'd27;
        rom[457][26] = -8'd4;
        rom[457][27] = 8'd9;
        rom[457][28] = -8'd5;
        rom[457][29] = -8'd3;
        rom[457][30] = -8'd76;
        rom[457][31] = 8'd13;
        rom[457][32] = -8'd7;
        rom[457][33] = -8'd28;
        rom[457][34] = 8'd20;
        rom[457][35] = 8'd2;
        rom[457][36] = -8'd34;
        rom[457][37] = -8'd36;
        rom[457][38] = -8'd5;
        rom[457][39] = -8'd22;
        rom[457][40] = 8'd13;
        rom[457][41] = 8'd41;
        rom[457][42] = -8'd14;
        rom[457][43] = -8'd9;
        rom[457][44] = -8'd39;
        rom[457][45] = -8'd11;
        rom[457][46] = -8'd37;
        rom[457][47] = 8'd30;
        rom[457][48] = 8'd42;
        rom[457][49] = -8'd21;
        rom[457][50] = -8'd6;
        rom[457][51] = 8'd23;
        rom[457][52] = -8'd10;
        rom[457][53] = 8'd3;
        rom[457][54] = 8'd7;
        rom[457][55] = -8'd10;
        rom[457][56] = -8'd21;
        rom[457][57] = 8'd32;
        rom[457][58] = 8'd39;
        rom[457][59] = -8'd27;
        rom[457][60] = -8'd20;
        rom[457][61] = 8'd11;
        rom[457][62] = 8'd36;
        rom[457][63] = 8'd0;
        rom[458][0] = 8'd10;
        rom[458][1] = -8'd22;
        rom[458][2] = -8'd13;
        rom[458][3] = 8'd21;
        rom[458][4] = -8'd41;
        rom[458][5] = -8'd4;
        rom[458][6] = -8'd35;
        rom[458][7] = -8'd5;
        rom[458][8] = 8'd22;
        rom[458][9] = 8'd3;
        rom[458][10] = 8'd22;
        rom[458][11] = -8'd20;
        rom[458][12] = -8'd2;
        rom[458][13] = 8'd11;
        rom[458][14] = -8'd63;
        rom[458][15] = 8'd49;
        rom[458][16] = -8'd10;
        rom[458][17] = -8'd7;
        rom[458][18] = -8'd36;
        rom[458][19] = -8'd23;
        rom[458][20] = -8'd13;
        rom[458][21] = -8'd32;
        rom[458][22] = -8'd12;
        rom[458][23] = -8'd49;
        rom[458][24] = 8'd10;
        rom[458][25] = 8'd11;
        rom[458][26] = -8'd11;
        rom[458][27] = 8'd21;
        rom[458][28] = 8'd41;
        rom[458][29] = 8'd22;
        rom[458][30] = 8'd10;
        rom[458][31] = 8'd21;
        rom[458][32] = 8'd13;
        rom[458][33] = 8'd5;
        rom[458][34] = -8'd8;
        rom[458][35] = 8'd5;
        rom[458][36] = -8'd23;
        rom[458][37] = 8'd38;
        rom[458][38] = -8'd30;
        rom[458][39] = -8'd43;
        rom[458][40] = -8'd7;
        rom[458][41] = -8'd22;
        rom[458][42] = 8'd0;
        rom[458][43] = 8'd2;
        rom[458][44] = 8'd8;
        rom[458][45] = 8'd0;
        rom[458][46] = 8'd21;
        rom[458][47] = 8'd10;
        rom[458][48] = -8'd3;
        rom[458][49] = -8'd18;
        rom[458][50] = 8'd0;
        rom[458][51] = -8'd16;
        rom[458][52] = -8'd3;
        rom[458][53] = -8'd37;
        rom[458][54] = -8'd7;
        rom[458][55] = -8'd12;
        rom[458][56] = 8'd5;
        rom[458][57] = -8'd34;
        rom[458][58] = 8'd13;
        rom[458][59] = 8'd36;
        rom[458][60] = 8'd4;
        rom[458][61] = -8'd48;
        rom[458][62] = 8'd36;
        rom[458][63] = -8'd3;
        rom[459][0] = -8'd45;
        rom[459][1] = -8'd11;
        rom[459][2] = 8'd6;
        rom[459][3] = -8'd49;
        rom[459][4] = 8'd47;
        rom[459][5] = -8'd1;
        rom[459][6] = -8'd14;
        rom[459][7] = -8'd50;
        rom[459][8] = -8'd41;
        rom[459][9] = -8'd4;
        rom[459][10] = 8'd17;
        rom[459][11] = -8'd42;
        rom[459][12] = -8'd26;
        rom[459][13] = -8'd45;
        rom[459][14] = 8'd27;
        rom[459][15] = 8'd0;
        rom[459][16] = -8'd6;
        rom[459][17] = -8'd23;
        rom[459][18] = -8'd64;
        rom[459][19] = 8'd12;
        rom[459][20] = -8'd5;
        rom[459][21] = -8'd26;
        rom[459][22] = 8'd14;
        rom[459][23] = -8'd36;
        rom[459][24] = -8'd14;
        rom[459][25] = 8'd10;
        rom[459][26] = 8'd25;
        rom[459][27] = 8'd7;
        rom[459][28] = 8'd11;
        rom[459][29] = -8'd13;
        rom[459][30] = 8'd26;
        rom[459][31] = -8'd28;
        rom[459][32] = -8'd22;
        rom[459][33] = -8'd15;
        rom[459][34] = -8'd3;
        rom[459][35] = -8'd6;
        rom[459][36] = -8'd10;
        rom[459][37] = 8'd6;
        rom[459][38] = -8'd23;
        rom[459][39] = -8'd5;
        rom[459][40] = -8'd32;
        rom[459][41] = 8'd40;
        rom[459][42] = 8'd22;
        rom[459][43] = 8'd18;
        rom[459][44] = -8'd16;
        rom[459][45] = -8'd38;
        rom[459][46] = 8'd8;
        rom[459][47] = 8'd13;
        rom[459][48] = -8'd17;
        rom[459][49] = -8'd23;
        rom[459][50] = -8'd57;
        rom[459][51] = 8'd4;
        rom[459][52] = 8'd51;
        rom[459][53] = -8'd54;
        rom[459][54] = -8'd14;
        rom[459][55] = -8'd35;
        rom[459][56] = 8'd0;
        rom[459][57] = -8'd35;
        rom[459][58] = -8'd11;
        rom[459][59] = -8'd29;
        rom[459][60] = -8'd13;
        rom[459][61] = -8'd13;
        rom[459][62] = 8'd34;
        rom[459][63] = -8'd35;
        rom[460][0] = -8'd111;
        rom[460][1] = -8'd55;
        rom[460][2] = -8'd61;
        rom[460][3] = 8'd22;
        rom[460][4] = 8'd25;
        rom[460][5] = -8'd4;
        rom[460][6] = 8'd14;
        rom[460][7] = 8'd55;
        rom[460][8] = 8'd26;
        rom[460][9] = 8'd5;
        rom[460][10] = 8'd15;
        rom[460][11] = -8'd15;
        rom[460][12] = -8'd9;
        rom[460][13] = -8'd84;
        rom[460][14] = 8'd15;
        rom[460][15] = 8'd23;
        rom[460][16] = 8'd29;
        rom[460][17] = -8'd16;
        rom[460][18] = 8'd11;
        rom[460][19] = -8'd49;
        rom[460][20] = -8'd4;
        rom[460][21] = 8'd36;
        rom[460][22] = -8'd20;
        rom[460][23] = -8'd34;
        rom[460][24] = 8'd5;
        rom[460][25] = 8'd9;
        rom[460][26] = -8'd4;
        rom[460][27] = 8'd33;
        rom[460][28] = 8'd5;
        rom[460][29] = -8'd3;
        rom[460][30] = 8'd21;
        rom[460][31] = -8'd20;
        rom[460][32] = 8'd13;
        rom[460][33] = -8'd37;
        rom[460][34] = 8'd16;
        rom[460][35] = 8'd20;
        rom[460][36] = -8'd15;
        rom[460][37] = -8'd4;
        rom[460][38] = 8'd8;
        rom[460][39] = 8'd2;
        rom[460][40] = -8'd49;
        rom[460][41] = -8'd3;
        rom[460][42] = -8'd17;
        rom[460][43] = 8'd1;
        rom[460][44] = 8'd0;
        rom[460][45] = 8'd11;
        rom[460][46] = 8'd17;
        rom[460][47] = 8'd9;
        rom[460][48] = -8'd26;
        rom[460][49] = 8'd4;
        rom[460][50] = 8'd34;
        rom[460][51] = 8'd20;
        rom[460][52] = -8'd48;
        rom[460][53] = -8'd10;
        rom[460][54] = 8'd7;
        rom[460][55] = -8'd15;
        rom[460][56] = -8'd57;
        rom[460][57] = -8'd6;
        rom[460][58] = 8'd13;
        rom[460][59] = 8'd8;
        rom[460][60] = 8'd0;
        rom[460][61] = 8'd16;
        rom[460][62] = -8'd4;
        rom[460][63] = 8'd3;
        rom[461][0] = 8'd5;
        rom[461][1] = 8'd18;
        rom[461][2] = 8'd1;
        rom[461][3] = 8'd15;
        rom[461][4] = 8'd0;
        rom[461][5] = 8'd41;
        rom[461][6] = -8'd12;
        rom[461][7] = 8'd10;
        rom[461][8] = -8'd1;
        rom[461][9] = 8'd14;
        rom[461][10] = 8'd7;
        rom[461][11] = -8'd41;
        rom[461][12] = -8'd46;
        rom[461][13] = -8'd38;
        rom[461][14] = -8'd37;
        rom[461][15] = 8'd17;
        rom[461][16] = -8'd46;
        rom[461][17] = -8'd42;
        rom[461][18] = -8'd7;
        rom[461][19] = -8'd1;
        rom[461][20] = -8'd13;
        rom[461][21] = -8'd10;
        rom[461][22] = -8'd25;
        rom[461][23] = 8'd11;
        rom[461][24] = 8'd19;
        rom[461][25] = 8'd18;
        rom[461][26] = 8'd18;
        rom[461][27] = 8'd52;
        rom[461][28] = -8'd8;
        rom[461][29] = 8'd20;
        rom[461][30] = -8'd32;
        rom[461][31] = 8'd3;
        rom[461][32] = -8'd15;
        rom[461][33] = 8'd14;
        rom[461][34] = -8'd13;
        rom[461][35] = -8'd29;
        rom[461][36] = -8'd17;
        rom[461][37] = -8'd10;
        rom[461][38] = -8'd3;
        rom[461][39] = 8'd3;
        rom[461][40] = 8'd28;
        rom[461][41] = 8'd13;
        rom[461][42] = -8'd17;
        rom[461][43] = 8'd15;
        rom[461][44] = 8'd10;
        rom[461][45] = 8'd18;
        rom[461][46] = -8'd20;
        rom[461][47] = -8'd18;
        rom[461][48] = 8'd31;
        rom[461][49] = -8'd23;
        rom[461][50] = 8'd5;
        rom[461][51] = -8'd26;
        rom[461][52] = 8'd11;
        rom[461][53] = -8'd12;
        rom[461][54] = -8'd25;
        rom[461][55] = -8'd14;
        rom[461][56] = -8'd9;
        rom[461][57] = -8'd47;
        rom[461][58] = 8'd25;
        rom[461][59] = 8'd7;
        rom[461][60] = 8'd10;
        rom[461][61] = -8'd42;
        rom[461][62] = 8'd42;
        rom[461][63] = -8'd21;
        rom[462][0] = -8'd4;
        rom[462][1] = -8'd24;
        rom[462][2] = 8'd10;
        rom[462][3] = -8'd26;
        rom[462][4] = 8'd5;
        rom[462][5] = -8'd42;
        rom[462][6] = 8'd8;
        rom[462][7] = -8'd59;
        rom[462][8] = -8'd6;
        rom[462][9] = -8'd69;
        rom[462][10] = -8'd16;
        rom[462][11] = -8'd42;
        rom[462][12] = -8'd7;
        rom[462][13] = -8'd6;
        rom[462][14] = -8'd1;
        rom[462][15] = -8'd6;
        rom[462][16] = -8'd32;
        rom[462][17] = 8'd27;
        rom[462][18] = -8'd5;
        rom[462][19] = 8'd27;
        rom[462][20] = -8'd2;
        rom[462][21] = -8'd29;
        rom[462][22] = 8'd37;
        rom[462][23] = -8'd21;
        rom[462][24] = 8'd12;
        rom[462][25] = -8'd11;
        rom[462][26] = -8'd16;
        rom[462][27] = -8'd38;
        rom[462][28] = -8'd18;
        rom[462][29] = -8'd23;
        rom[462][30] = 8'd1;
        rom[462][31] = 8'd2;
        rom[462][32] = 8'd23;
        rom[462][33] = -8'd27;
        rom[462][34] = -8'd1;
        rom[462][35] = 8'd10;
        rom[462][36] = -8'd4;
        rom[462][37] = 8'd18;
        rom[462][38] = -8'd5;
        rom[462][39] = 8'd28;
        rom[462][40] = 8'd9;
        rom[462][41] = -8'd22;
        rom[462][42] = 8'd11;
        rom[462][43] = 8'd2;
        rom[462][44] = 8'd17;
        rom[462][45] = -8'd24;
        rom[462][46] = -8'd25;
        rom[462][47] = 8'd20;
        rom[462][48] = -8'd4;
        rom[462][49] = -8'd12;
        rom[462][50] = -8'd16;
        rom[462][51] = 8'd8;
        rom[462][52] = -8'd30;
        rom[462][53] = -8'd21;
        rom[462][54] = 8'd38;
        rom[462][55] = 8'd18;
        rom[462][56] = -8'd10;
        rom[462][57] = -8'd1;
        rom[462][58] = 8'd19;
        rom[462][59] = -8'd42;
        rom[462][60] = 8'd19;
        rom[462][61] = 8'd2;
        rom[462][62] = 8'd29;
        rom[462][63] = 8'd23;
        rom[463][0] = 8'd13;
        rom[463][1] = -8'd17;
        rom[463][2] = 8'd52;
        rom[463][3] = -8'd21;
        rom[463][4] = 8'd40;
        rom[463][5] = 8'd16;
        rom[463][6] = -8'd14;
        rom[463][7] = -8'd30;
        rom[463][8] = 8'd13;
        rom[463][9] = 8'd0;
        rom[463][10] = -8'd58;
        rom[463][11] = 8'd0;
        rom[463][12] = 8'd37;
        rom[463][13] = -8'd8;
        rom[463][14] = -8'd15;
        rom[463][15] = 8'd8;
        rom[463][16] = -8'd15;
        rom[463][17] = 8'd28;
        rom[463][18] = -8'd2;
        rom[463][19] = -8'd22;
        rom[463][20] = -8'd13;
        rom[463][21] = -8'd48;
        rom[463][22] = -8'd4;
        rom[463][23] = -8'd1;
        rom[463][24] = -8'd25;
        rom[463][25] = -8'd40;
        rom[463][26] = -8'd21;
        rom[463][27] = 8'd17;
        rom[463][28] = 8'd7;
        rom[463][29] = -8'd12;
        rom[463][30] = -8'd7;
        rom[463][31] = -8'd9;
        rom[463][32] = -8'd4;
        rom[463][33] = -8'd13;
        rom[463][34] = -8'd12;
        rom[463][35] = 8'd9;
        rom[463][36] = -8'd22;
        rom[463][37] = -8'd99;
        rom[463][38] = -8'd20;
        rom[463][39] = 8'd7;
        rom[463][40] = 8'd16;
        rom[463][41] = 8'd8;
        rom[463][42] = 8'd2;
        rom[463][43] = 8'd18;
        rom[463][44] = 8'd38;
        rom[463][45] = -8'd25;
        rom[463][46] = 8'd2;
        rom[463][47] = 8'd9;
        rom[463][48] = 8'd16;
        rom[463][49] = -8'd1;
        rom[463][50] = 8'd17;
        rom[463][51] = 8'd18;
        rom[463][52] = 8'd0;
        rom[463][53] = 8'd27;
        rom[463][54] = 8'd10;
        rom[463][55] = -8'd21;
        rom[463][56] = -8'd21;
        rom[463][57] = -8'd14;
        rom[463][58] = -8'd34;
        rom[463][59] = 8'd11;
        rom[463][60] = -8'd2;
        rom[463][61] = -8'd30;
        rom[463][62] = -8'd11;
        rom[463][63] = 8'd10;
        rom[464][0] = -8'd6;
        rom[464][1] = -8'd4;
        rom[464][2] = -8'd9;
        rom[464][3] = -8'd9;
        rom[464][4] = -8'd3;
        rom[464][5] = 8'd9;
        rom[464][6] = 8'd3;
        rom[464][7] = 8'd9;
        rom[464][8] = 8'd4;
        rom[464][9] = 8'd4;
        rom[464][10] = 8'd1;
        rom[464][11] = 8'd2;
        rom[464][12] = 8'd0;
        rom[464][13] = -8'd2;
        rom[464][14] = -8'd7;
        rom[464][15] = -8'd2;
        rom[464][16] = -8'd7;
        rom[464][17] = -8'd1;
        rom[464][18] = -8'd7;
        rom[464][19] = -8'd5;
        rom[464][20] = -8'd6;
        rom[464][21] = -8'd4;
        rom[464][22] = 8'd4;
        rom[464][23] = -8'd1;
        rom[464][24] = 8'd5;
        rom[464][25] = 8'd1;
        rom[464][26] = -8'd1;
        rom[464][27] = -8'd7;
        rom[464][28] = -8'd5;
        rom[464][29] = 8'd2;
        rom[464][30] = 8'd0;
        rom[464][31] = 8'd6;
        rom[464][32] = -8'd5;
        rom[464][33] = 8'd5;
        rom[464][34] = -8'd5;
        rom[464][35] = 8'd1;
        rom[464][36] = -8'd8;
        rom[464][37] = -8'd3;
        rom[464][38] = -8'd4;
        rom[464][39] = -8'd2;
        rom[464][40] = -8'd4;
        rom[464][41] = 8'd0;
        rom[464][42] = 8'd9;
        rom[464][43] = 8'd4;
        rom[464][44] = 8'd2;
        rom[464][45] = -8'd9;
        rom[464][46] = -8'd2;
        rom[464][47] = 8'd2;
        rom[464][48] = -8'd8;
        rom[464][49] = -8'd8;
        rom[464][50] = -8'd3;
        rom[464][51] = -8'd5;
        rom[464][52] = -8'd9;
        rom[464][53] = 8'd6;
        rom[464][54] = 8'd8;
        rom[464][55] = 8'd6;
        rom[464][56] = 8'd4;
        rom[464][57] = -8'd7;
        rom[464][58] = 8'd0;
        rom[464][59] = -8'd4;
        rom[464][60] = -8'd5;
        rom[464][61] = 8'd8;
        rom[464][62] = -8'd8;
        rom[464][63] = 8'd7;
        rom[465][0] = 8'd11;
        rom[465][1] = 8'd0;
        rom[465][2] = -8'd30;
        rom[465][3] = 8'd22;
        rom[465][4] = -8'd15;
        rom[465][5] = 8'd5;
        rom[465][6] = -8'd9;
        rom[465][7] = -8'd22;
        rom[465][8] = -8'd24;
        rom[465][9] = -8'd12;
        rom[465][10] = -8'd62;
        rom[465][11] = 8'd6;
        rom[465][12] = -8'd10;
        rom[465][13] = 8'd35;
        rom[465][14] = -8'd8;
        rom[465][15] = -8'd16;
        rom[465][16] = 8'd4;
        rom[465][17] = 8'd17;
        rom[465][18] = 8'd17;
        rom[465][19] = 8'd6;
        rom[465][20] = -8'd9;
        rom[465][21] = -8'd16;
        rom[465][22] = -8'd25;
        rom[465][23] = -8'd18;
        rom[465][24] = 8'd21;
        rom[465][25] = 8'd22;
        rom[465][26] = -8'd35;
        rom[465][27] = -8'd43;
        rom[465][28] = -8'd32;
        rom[465][29] = -8'd66;
        rom[465][30] = -8'd4;
        rom[465][31] = 8'd25;
        rom[465][32] = -8'd2;
        rom[465][33] = 8'd11;
        rom[465][34] = -8'd24;
        rom[465][35] = -8'd5;
        rom[465][36] = 8'd43;
        rom[465][37] = 8'd3;
        rom[465][38] = -8'd43;
        rom[465][39] = -8'd8;
        rom[465][40] = -8'd16;
        rom[465][41] = -8'd16;
        rom[465][42] = -8'd29;
        rom[465][43] = -8'd2;
        rom[465][44] = 8'd28;
        rom[465][45] = 8'd45;
        rom[465][46] = -8'd4;
        rom[465][47] = -8'd17;
        rom[465][48] = 8'd13;
        rom[465][49] = 8'd10;
        rom[465][50] = -8'd9;
        rom[465][51] = -8'd7;
        rom[465][52] = 8'd26;
        rom[465][53] = -8'd20;
        rom[465][54] = 8'd10;
        rom[465][55] = 8'd0;
        rom[465][56] = -8'd6;
        rom[465][57] = -8'd28;
        rom[465][58] = -8'd33;
        rom[465][59] = 8'd21;
        rom[465][60] = 8'd28;
        rom[465][61] = 8'd62;
        rom[465][62] = -8'd1;
        rom[465][63] = -8'd33;
        rom[466][0] = 8'd59;
        rom[466][1] = -8'd24;
        rom[466][2] = 8'd20;
        rom[466][3] = -8'd39;
        rom[466][4] = 8'd10;
        rom[466][5] = 8'd19;
        rom[466][6] = 8'd20;
        rom[466][7] = 8'd7;
        rom[466][8] = 8'd18;
        rom[466][9] = -8'd22;
        rom[466][10] = -8'd23;
        rom[466][11] = 8'd11;
        rom[466][12] = -8'd54;
        rom[466][13] = -8'd14;
        rom[466][14] = -8'd1;
        rom[466][15] = -8'd16;
        rom[466][16] = -8'd70;
        rom[466][17] = -8'd87;
        rom[466][18] = 8'd1;
        rom[466][19] = 8'd8;
        rom[466][20] = -8'd4;
        rom[466][21] = -8'd9;
        rom[466][22] = -8'd14;
        rom[466][23] = 8'd33;
        rom[466][24] = -8'd1;
        rom[466][25] = -8'd28;
        rom[466][26] = -8'd34;
        rom[466][27] = -8'd19;
        rom[466][28] = -8'd29;
        rom[466][29] = -8'd24;
        rom[466][30] = -8'd35;
        rom[466][31] = -8'd13;
        rom[466][32] = 8'd14;
        rom[466][33] = -8'd14;
        rom[466][34] = 8'd13;
        rom[466][35] = -8'd2;
        rom[466][36] = 8'd2;
        rom[466][37] = -8'd45;
        rom[466][38] = -8'd51;
        rom[466][39] = 8'd22;
        rom[466][40] = -8'd39;
        rom[466][41] = 8'd14;
        rom[466][42] = -8'd2;
        rom[466][43] = -8'd2;
        rom[466][44] = 8'd15;
        rom[466][45] = -8'd54;
        rom[466][46] = -8'd34;
        rom[466][47] = -8'd74;
        rom[466][48] = -8'd19;
        rom[466][49] = -8'd13;
        rom[466][50] = -8'd12;
        rom[466][51] = -8'd20;
        rom[466][52] = -8'd17;
        rom[466][53] = 8'd2;
        rom[466][54] = 8'd24;
        rom[466][55] = 8'd9;
        rom[466][56] = 8'd3;
        rom[466][57] = -8'd10;
        rom[466][58] = -8'd18;
        rom[466][59] = -8'd3;
        rom[466][60] = -8'd20;
        rom[466][61] = 8'd4;
        rom[466][62] = 8'd9;
        rom[466][63] = 8'd37;
        rom[467][0] = 8'd26;
        rom[467][1] = -8'd14;
        rom[467][2] = 8'd4;
        rom[467][3] = -8'd16;
        rom[467][4] = -8'd38;
        rom[467][5] = -8'd12;
        rom[467][6] = -8'd22;
        rom[467][7] = 8'd30;
        rom[467][8] = -8'd26;
        rom[467][9] = -8'd45;
        rom[467][10] = 8'd1;
        rom[467][11] = -8'd33;
        rom[467][12] = 8'd0;
        rom[467][13] = 8'd30;
        rom[467][14] = 8'd2;
        rom[467][15] = 8'd45;
        rom[467][16] = 8'd26;
        rom[467][17] = 8'd5;
        rom[467][18] = -8'd20;
        rom[467][19] = 8'd5;
        rom[467][20] = 8'd5;
        rom[467][21] = -8'd24;
        rom[467][22] = -8'd15;
        rom[467][23] = 8'd2;
        rom[467][24] = 8'd17;
        rom[467][25] = 8'd8;
        rom[467][26] = -8'd8;
        rom[467][27] = 8'd6;
        rom[467][28] = -8'd18;
        rom[467][29] = 8'd26;
        rom[467][30] = 8'd7;
        rom[467][31] = -8'd64;
        rom[467][32] = 8'd11;
        rom[467][33] = 8'd2;
        rom[467][34] = 8'd13;
        rom[467][35] = -8'd73;
        rom[467][36] = 8'd34;
        rom[467][37] = -8'd51;
        rom[467][38] = -8'd20;
        rom[467][39] = -8'd13;
        rom[467][40] = 8'd18;
        rom[467][41] = -8'd28;
        rom[467][42] = 8'd18;
        rom[467][43] = -8'd8;
        rom[467][44] = 8'd15;
        rom[467][45] = -8'd18;
        rom[467][46] = 8'd7;
        rom[467][47] = -8'd10;
        rom[467][48] = 8'd18;
        rom[467][49] = -8'd28;
        rom[467][50] = -8'd15;
        rom[467][51] = 8'd26;
        rom[467][52] = 8'd15;
        rom[467][53] = 8'd3;
        rom[467][54] = -8'd22;
        rom[467][55] = -8'd15;
        rom[467][56] = -8'd20;
        rom[467][57] = 8'd20;
        rom[467][58] = -8'd23;
        rom[467][59] = 8'd7;
        rom[467][60] = -8'd42;
        rom[467][61] = 8'd0;
        rom[467][62] = 8'd31;
        rom[467][63] = -8'd27;
        rom[468][0] = -8'd35;
        rom[468][1] = -8'd10;
        rom[468][2] = -8'd22;
        rom[468][3] = 8'd1;
        rom[468][4] = -8'd106;
        rom[468][5] = 8'd15;
        rom[468][6] = -8'd20;
        rom[468][7] = -8'd3;
        rom[468][8] = -8'd16;
        rom[468][9] = -8'd42;
        rom[468][10] = 8'd4;
        rom[468][11] = -8'd1;
        rom[468][12] = 8'd5;
        rom[468][13] = -8'd15;
        rom[468][14] = -8'd58;
        rom[468][15] = -8'd9;
        rom[468][16] = -8'd13;
        rom[468][17] = -8'd23;
        rom[468][18] = -8'd20;
        rom[468][19] = 8'd6;
        rom[468][20] = 8'd1;
        rom[468][21] = 8'd1;
        rom[468][22] = -8'd59;
        rom[468][23] = -8'd70;
        rom[468][24] = 8'd23;
        rom[468][25] = -8'd5;
        rom[468][26] = 8'd4;
        rom[468][27] = -8'd4;
        rom[468][28] = -8'd21;
        rom[468][29] = -8'd21;
        rom[468][30] = -8'd41;
        rom[468][31] = -8'd31;
        rom[468][32] = 8'd0;
        rom[468][33] = -8'd6;
        rom[468][34] = 8'd11;
        rom[468][35] = -8'd65;
        rom[468][36] = -8'd12;
        rom[468][37] = -8'd19;
        rom[468][38] = 8'd10;
        rom[468][39] = -8'd1;
        rom[468][40] = 8'd4;
        rom[468][41] = -8'd35;
        rom[468][42] = 8'd44;
        rom[468][43] = -8'd2;
        rom[468][44] = 8'd13;
        rom[468][45] = -8'd44;
        rom[468][46] = -8'd6;
        rom[468][47] = -8'd2;
        rom[468][48] = -8'd54;
        rom[468][49] = 8'd12;
        rom[468][50] = -8'd49;
        rom[468][51] = 8'd20;
        rom[468][52] = 8'd6;
        rom[468][53] = -8'd39;
        rom[468][54] = -8'd22;
        rom[468][55] = 8'd16;
        rom[468][56] = 8'd10;
        rom[468][57] = 8'd6;
        rom[468][58] = -8'd9;
        rom[468][59] = -8'd26;
        rom[468][60] = 8'd2;
        rom[468][61] = -8'd12;
        rom[468][62] = -8'd1;
        rom[468][63] = -8'd19;
        rom[469][0] = 8'd7;
        rom[469][1] = -8'd4;
        rom[469][2] = -8'd2;
        rom[469][3] = -8'd1;
        rom[469][4] = 8'd7;
        rom[469][5] = -8'd4;
        rom[469][6] = 8'd3;
        rom[469][7] = -8'd3;
        rom[469][8] = 8'd7;
        rom[469][9] = -8'd1;
        rom[469][10] = -8'd5;
        rom[469][11] = -8'd9;
        rom[469][12] = -8'd4;
        rom[469][13] = -8'd1;
        rom[469][14] = 8'd5;
        rom[469][15] = -8'd6;
        rom[469][16] = 8'd12;
        rom[469][17] = 8'd4;
        rom[469][18] = 8'd6;
        rom[469][19] = -8'd4;
        rom[469][20] = 8'd7;
        rom[469][21] = 8'd10;
        rom[469][22] = -8'd6;
        rom[469][23] = 8'd3;
        rom[469][24] = 8'd5;
        rom[469][25] = -8'd8;
        rom[469][26] = -8'd7;
        rom[469][27] = 8'd4;
        rom[469][28] = 8'd0;
        rom[469][29] = -8'd3;
        rom[469][30] = -8'd3;
        rom[469][31] = 8'd4;
        rom[469][32] = -8'd1;
        rom[469][33] = -8'd4;
        rom[469][34] = -8'd7;
        rom[469][35] = 8'd0;
        rom[469][36] = -8'd6;
        rom[469][37] = -8'd9;
        rom[469][38] = 8'd2;
        rom[469][39] = 8'd2;
        rom[469][40] = -8'd8;
        rom[469][41] = -8'd2;
        rom[469][42] = -8'd11;
        rom[469][43] = 8'd0;
        rom[469][44] = 8'd7;
        rom[469][45] = 8'd6;
        rom[469][46] = -8'd4;
        rom[469][47] = 8'd11;
        rom[469][48] = -8'd5;
        rom[469][49] = 8'd2;
        rom[469][50] = 8'd7;
        rom[469][51] = 8'd5;
        rom[469][52] = -8'd9;
        rom[469][53] = 8'd1;
        rom[469][54] = -8'd9;
        rom[469][55] = 8'd1;
        rom[469][56] = 8'd6;
        rom[469][57] = -8'd4;
        rom[469][58] = -8'd1;
        rom[469][59] = -8'd4;
        rom[469][60] = 8'd1;
        rom[469][61] = 8'd2;
        rom[469][62] = -8'd4;
        rom[469][63] = 8'd5;
        rom[470][0] = -8'd69;
        rom[470][1] = 8'd26;
        rom[470][2] = -8'd5;
        rom[470][3] = 8'd27;
        rom[470][4] = -8'd12;
        rom[470][5] = -8'd4;
        rom[470][6] = 8'd23;
        rom[470][7] = -8'd63;
        rom[470][8] = 8'd13;
        rom[470][9] = 8'd14;
        rom[470][10] = 8'd22;
        rom[470][11] = -8'd13;
        rom[470][12] = -8'd63;
        rom[470][13] = -8'd15;
        rom[470][14] = -8'd1;
        rom[470][15] = -8'd18;
        rom[470][16] = 8'd31;
        rom[470][17] = 8'd15;
        rom[470][18] = -8'd32;
        rom[470][19] = 8'd15;
        rom[470][20] = -8'd1;
        rom[470][21] = -8'd19;
        rom[470][22] = -8'd37;
        rom[470][23] = 8'd13;
        rom[470][24] = -8'd31;
        rom[470][25] = 8'd22;
        rom[470][26] = 8'd34;
        rom[470][27] = 8'd20;
        rom[470][28] = -8'd3;
        rom[470][29] = 8'd21;
        rom[470][30] = -8'd36;
        rom[470][31] = 8'd2;
        rom[470][32] = -8'd9;
        rom[470][33] = 8'd23;
        rom[470][34] = 8'd12;
        rom[470][35] = -8'd20;
        rom[470][36] = -8'd37;
        rom[470][37] = 8'd9;
        rom[470][38] = 8'd13;
        rom[470][39] = 8'd10;
        rom[470][40] = 8'd32;
        rom[470][41] = 8'd0;
        rom[470][42] = -8'd19;
        rom[470][43] = -8'd25;
        rom[470][44] = -8'd24;
        rom[470][45] = -8'd7;
        rom[470][46] = -8'd24;
        rom[470][47] = -8'd39;
        rom[470][48] = -8'd45;
        rom[470][49] = -8'd8;
        rom[470][50] = -8'd10;
        rom[470][51] = -8'd12;
        rom[470][52] = 8'd18;
        rom[470][53] = 8'd5;
        rom[470][54] = 8'd1;
        rom[470][55] = -8'd8;
        rom[470][56] = -8'd35;
        rom[470][57] = -8'd1;
        rom[470][58] = 8'd10;
        rom[470][59] = 8'd17;
        rom[470][60] = 8'd11;
        rom[470][61] = 8'd14;
        rom[470][62] = -8'd39;
        rom[470][63] = 8'd27;
        rom[471][0] = -8'd21;
        rom[471][1] = 8'd10;
        rom[471][2] = 8'd13;
        rom[471][3] = 8'd3;
        rom[471][4] = 8'd45;
        rom[471][5] = 8'd1;
        rom[471][6] = 8'd3;
        rom[471][7] = -8'd2;
        rom[471][8] = -8'd17;
        rom[471][9] = 8'd12;
        rom[471][10] = 8'd30;
        rom[471][11] = -8'd10;
        rom[471][12] = 8'd33;
        rom[471][13] = -8'd7;
        rom[471][14] = -8'd44;
        rom[471][15] = -8'd18;
        rom[471][16] = -8'd38;
        rom[471][17] = -8'd29;
        rom[471][18] = -8'd13;
        rom[471][19] = -8'd20;
        rom[471][20] = -8'd10;
        rom[471][21] = 8'd18;
        rom[471][22] = -8'd20;
        rom[471][23] = -8'd12;
        rom[471][24] = -8'd26;
        rom[471][25] = -8'd23;
        rom[471][26] = -8'd46;
        rom[471][27] = -8'd3;
        rom[471][28] = 8'd51;
        rom[471][29] = -8'd3;
        rom[471][30] = 8'd20;
        rom[471][31] = -8'd46;
        rom[471][32] = 8'd33;
        rom[471][33] = -8'd26;
        rom[471][34] = 8'd32;
        rom[471][35] = -8'd5;
        rom[471][36] = -8'd22;
        rom[471][37] = -8'd8;
        rom[471][38] = 8'd8;
        rom[471][39] = -8'd6;
        rom[471][40] = -8'd28;
        rom[471][41] = -8'd12;
        rom[471][42] = 8'd9;
        rom[471][43] = 8'd13;
        rom[471][44] = -8'd18;
        rom[471][45] = -8'd29;
        rom[471][46] = 8'd38;
        rom[471][47] = 8'd28;
        rom[471][48] = -8'd69;
        rom[471][49] = 8'd10;
        rom[471][50] = -8'd27;
        rom[471][51] = -8'd20;
        rom[471][52] = 8'd22;
        rom[471][53] = 8'd15;
        rom[471][54] = 8'd21;
        rom[471][55] = 8'd23;
        rom[471][56] = 8'd3;
        rom[471][57] = 8'd4;
        rom[471][58] = -8'd9;
        rom[471][59] = 8'd24;
        rom[471][60] = 8'd8;
        rom[471][61] = -8'd7;
        rom[471][62] = -8'd54;
        rom[471][63] = -8'd34;
        rom[472][0] = -8'd36;
        rom[472][1] = -8'd42;
        rom[472][2] = 8'd21;
        rom[472][3] = 8'd55;
        rom[472][4] = 8'd57;
        rom[472][5] = -8'd25;
        rom[472][6] = 8'd49;
        rom[472][7] = 8'd13;
        rom[472][8] = -8'd47;
        rom[472][9] = 8'd33;
        rom[472][10] = -8'd15;
        rom[472][11] = 8'd20;
        rom[472][12] = 8'd17;
        rom[472][13] = 8'd15;
        rom[472][14] = -8'd26;
        rom[472][15] = -8'd3;
        rom[472][16] = 8'd14;
        rom[472][17] = -8'd3;
        rom[472][18] = 8'd9;
        rom[472][19] = 8'd24;
        rom[472][20] = -8'd9;
        rom[472][21] = 8'd5;
        rom[472][22] = -8'd45;
        rom[472][23] = 8'd9;
        rom[472][24] = 8'd19;
        rom[472][25] = -8'd81;
        rom[472][26] = 8'd21;
        rom[472][27] = -8'd2;
        rom[472][28] = 8'd40;
        rom[472][29] = -8'd25;
        rom[472][30] = 8'd29;
        rom[472][31] = -8'd21;
        rom[472][32] = 8'd37;
        rom[472][33] = 8'd33;
        rom[472][34] = -8'd38;
        rom[472][35] = 8'd12;
        rom[472][36] = -8'd10;
        rom[472][37] = 8'd23;
        rom[472][38] = -8'd29;
        rom[472][39] = 8'd37;
        rom[472][40] = 8'd24;
        rom[472][41] = -8'd18;
        rom[472][42] = 8'd23;
        rom[472][43] = -8'd4;
        rom[472][44] = -8'd37;
        rom[472][45] = -8'd1;
        rom[472][46] = 8'd5;
        rom[472][47] = 8'd8;
        rom[472][48] = -8'd10;
        rom[472][49] = 8'd9;
        rom[472][50] = 8'd7;
        rom[472][51] = -8'd21;
        rom[472][52] = 8'd13;
        rom[472][53] = 8'd4;
        rom[472][54] = 8'd23;
        rom[472][55] = -8'd34;
        rom[472][56] = 8'd2;
        rom[472][57] = -8'd12;
        rom[472][58] = -8'd41;
        rom[472][59] = -8'd16;
        rom[472][60] = 8'd3;
        rom[472][61] = 8'd19;
        rom[472][62] = 8'd16;
        rom[472][63] = -8'd12;
        rom[473][0] = 8'd10;
        rom[473][1] = -8'd6;
        rom[473][2] = -8'd29;
        rom[473][3] = -8'd22;
        rom[473][4] = -8'd39;
        rom[473][5] = 8'd25;
        rom[473][6] = 8'd3;
        rom[473][7] = 8'd8;
        rom[473][8] = -8'd41;
        rom[473][9] = -8'd23;
        rom[473][10] = -8'd34;
        rom[473][11] = 8'd23;
        rom[473][12] = -8'd53;
        rom[473][13] = -8'd43;
        rom[473][14] = -8'd4;
        rom[473][15] = -8'd3;
        rom[473][16] = -8'd6;
        rom[473][17] = -8'd16;
        rom[473][18] = 8'd5;
        rom[473][19] = 8'd19;
        rom[473][20] = -8'd6;
        rom[473][21] = 8'd11;
        rom[473][22] = -8'd2;
        rom[473][23] = 8'd44;
        rom[473][24] = 8'd20;
        rom[473][25] = -8'd16;
        rom[473][26] = 8'd29;
        rom[473][27] = -8'd38;
        rom[473][28] = -8'd3;
        rom[473][29] = -8'd10;
        rom[473][30] = -8'd38;
        rom[473][31] = 8'd1;
        rom[473][32] = 8'd7;
        rom[473][33] = -8'd20;
        rom[473][34] = 8'd25;
        rom[473][35] = -8'd18;
        rom[473][36] = -8'd10;
        rom[473][37] = -8'd14;
        rom[473][38] = -8'd8;
        rom[473][39] = 8'd4;
        rom[473][40] = -8'd19;
        rom[473][41] = -8'd17;
        rom[473][42] = -8'd15;
        rom[473][43] = -8'd53;
        rom[473][44] = -8'd40;
        rom[473][45] = -8'd13;
        rom[473][46] = -8'd14;
        rom[473][47] = 8'd9;
        rom[473][48] = -8'd54;
        rom[473][49] = -8'd18;
        rom[473][50] = -8'd76;
        rom[473][51] = -8'd23;
        rom[473][52] = -8'd22;
        rom[473][53] = -8'd46;
        rom[473][54] = -8'd23;
        rom[473][55] = -8'd18;
        rom[473][56] = -8'd32;
        rom[473][57] = -8'd28;
        rom[473][58] = 8'd19;
        rom[473][59] = 8'd6;
        rom[473][60] = -8'd1;
        rom[473][61] = -8'd12;
        rom[473][62] = 8'd14;
        rom[473][63] = 8'd31;
        rom[474][0] = 8'd10;
        rom[474][1] = -8'd17;
        rom[474][2] = -8'd26;
        rom[474][3] = -8'd7;
        rom[474][4] = 8'd19;
        rom[474][5] = 8'd0;
        rom[474][6] = 8'd24;
        rom[474][7] = -8'd61;
        rom[474][8] = 8'd17;
        rom[474][9] = 8'd8;
        rom[474][10] = 8'd47;
        rom[474][11] = -8'd36;
        rom[474][12] = 8'd1;
        rom[474][13] = -8'd10;
        rom[474][14] = 8'd27;
        rom[474][15] = -8'd34;
        rom[474][16] = -8'd22;
        rom[474][17] = 8'd16;
        rom[474][18] = 8'd21;
        rom[474][19] = -8'd30;
        rom[474][20] = -8'd4;
        rom[474][21] = 8'd30;
        rom[474][22] = 8'd2;
        rom[474][23] = -8'd13;
        rom[474][24] = 8'd8;
        rom[474][25] = -8'd8;
        rom[474][26] = -8'd5;
        rom[474][27] = -8'd23;
        rom[474][28] = -8'd12;
        rom[474][29] = -8'd11;
        rom[474][30] = 8'd40;
        rom[474][31] = -8'd25;
        rom[474][32] = 8'd16;
        rom[474][33] = -8'd19;
        rom[474][34] = 8'd24;
        rom[474][35] = -8'd9;
        rom[474][36] = 8'd24;
        rom[474][37] = -8'd11;
        rom[474][38] = 8'd9;
        rom[474][39] = 8'd11;
        rom[474][40] = -8'd19;
        rom[474][41] = 8'd15;
        rom[474][42] = -8'd22;
        rom[474][43] = -8'd4;
        rom[474][44] = -8'd11;
        rom[474][45] = -8'd25;
        rom[474][46] = -8'd46;
        rom[474][47] = 8'd33;
        rom[474][48] = -8'd13;
        rom[474][49] = 8'd14;
        rom[474][50] = -8'd29;
        rom[474][51] = -8'd25;
        rom[474][52] = -8'd19;
        rom[474][53] = 8'd17;
        rom[474][54] = -8'd80;
        rom[474][55] = 8'd23;
        rom[474][56] = -8'd16;
        rom[474][57] = 8'd0;
        rom[474][58] = -8'd26;
        rom[474][59] = -8'd18;
        rom[474][60] = 8'd52;
        rom[474][61] = 8'd35;
        rom[474][62] = -8'd11;
        rom[474][63] = -8'd21;
        rom[475][0] = -8'd14;
        rom[475][1] = 8'd46;
        rom[475][2] = 8'd7;
        rom[475][3] = 8'd9;
        rom[475][4] = -8'd10;
        rom[475][5] = 8'd49;
        rom[475][6] = 8'd25;
        rom[475][7] = -8'd19;
        rom[475][8] = 8'd23;
        rom[475][9] = -8'd12;
        rom[475][10] = 8'd9;
        rom[475][11] = 8'd10;
        rom[475][12] = -8'd29;
        rom[475][13] = -8'd12;
        rom[475][14] = -8'd9;
        rom[475][15] = 8'd17;
        rom[475][16] = -8'd89;
        rom[475][17] = -8'd23;
        rom[475][18] = 8'd3;
        rom[475][19] = 8'd23;
        rom[475][20] = -8'd4;
        rom[475][21] = 8'd13;
        rom[475][22] = -8'd18;
        rom[475][23] = -8'd2;
        rom[475][24] = 8'd15;
        rom[475][25] = 8'd6;
        rom[475][26] = 8'd25;
        rom[475][27] = -8'd32;
        rom[475][28] = -8'd13;
        rom[475][29] = 8'd12;
        rom[475][30] = -8'd30;
        rom[475][31] = 8'd7;
        rom[475][32] = -8'd9;
        rom[475][33] = -8'd9;
        rom[475][34] = 8'd5;
        rom[475][35] = -8'd4;
        rom[475][36] = -8'd9;
        rom[475][37] = -8'd83;
        rom[475][38] = -8'd15;
        rom[475][39] = 8'd1;
        rom[475][40] = 8'd1;
        rom[475][41] = -8'd11;
        rom[475][42] = 8'd10;
        rom[475][43] = -8'd25;
        rom[475][44] = 8'd12;
        rom[475][45] = 8'd20;
        rom[475][46] = 8'd13;
        rom[475][47] = -8'd18;
        rom[475][48] = 8'd19;
        rom[475][49] = -8'd5;
        rom[475][50] = -8'd12;
        rom[475][51] = 8'd5;
        rom[475][52] = -8'd14;
        rom[475][53] = -8'd4;
        rom[475][54] = 8'd1;
        rom[475][55] = -8'd57;
        rom[475][56] = 8'd16;
        rom[475][57] = -8'd35;
        rom[475][58] = 8'd3;
        rom[475][59] = 8'd23;
        rom[475][60] = -8'd12;
        rom[475][61] = 8'd4;
        rom[475][62] = 8'd19;
        rom[475][63] = -8'd21;
        rom[476][0] = -8'd25;
        rom[476][1] = 8'd30;
        rom[476][2] = 8'd8;
        rom[476][3] = 8'd5;
        rom[476][4] = 8'd17;
        rom[476][5] = -8'd51;
        rom[476][6] = -8'd42;
        rom[476][7] = 8'd40;
        rom[476][8] = -8'd10;
        rom[476][9] = 8'd19;
        rom[476][10] = 8'd15;
        rom[476][11] = -8'd17;
        rom[476][12] = -8'd23;
        rom[476][13] = 8'd5;
        rom[476][14] = -8'd40;
        rom[476][15] = -8'd1;
        rom[476][16] = 8'd24;
        rom[476][17] = 8'd1;
        rom[476][18] = -8'd35;
        rom[476][19] = -8'd41;
        rom[476][20] = -8'd13;
        rom[476][21] = 8'd5;
        rom[476][22] = 8'd14;
        rom[476][23] = 8'd4;
        rom[476][24] = -8'd29;
        rom[476][25] = 8'd5;
        rom[476][26] = -8'd43;
        rom[476][27] = -8'd32;
        rom[476][28] = -8'd25;
        rom[476][29] = 8'd15;
        rom[476][30] = 8'd8;
        rom[476][31] = 8'd12;
        rom[476][32] = -8'd22;
        rom[476][33] = -8'd5;
        rom[476][34] = -8'd9;
        rom[476][35] = 8'd3;
        rom[476][36] = 8'd21;
        rom[476][37] = -8'd20;
        rom[476][38] = -8'd10;
        rom[476][39] = -8'd10;
        rom[476][40] = -8'd51;
        rom[476][41] = -8'd51;
        rom[476][42] = -8'd29;
        rom[476][43] = 8'd30;
        rom[476][44] = 8'd10;
        rom[476][45] = 8'd42;
        rom[476][46] = -8'd4;
        rom[476][47] = 8'd21;
        rom[476][48] = 8'd13;
        rom[476][49] = -8'd2;
        rom[476][50] = -8'd3;
        rom[476][51] = -8'd19;
        rom[476][52] = -8'd7;
        rom[476][53] = 8'd4;
        rom[476][54] = -8'd15;
        rom[476][55] = 8'd32;
        rom[476][56] = 8'd16;
        rom[476][57] = -8'd29;
        rom[476][58] = -8'd16;
        rom[476][59] = 8'd16;
        rom[476][60] = -8'd57;
        rom[476][61] = -8'd16;
        rom[476][62] = 8'd35;
        rom[476][63] = 8'd2;
        rom[477][0] = 8'd40;
        rom[477][1] = -8'd22;
        rom[477][2] = 8'd24;
        rom[477][3] = 8'd5;
        rom[477][4] = -8'd61;
        rom[477][5] = -8'd11;
        rom[477][6] = 8'd15;
        rom[477][7] = 8'd44;
        rom[477][8] = 8'd11;
        rom[477][9] = -8'd12;
        rom[477][10] = 8'd38;
        rom[477][11] = -8'd29;
        rom[477][12] = -8'd19;
        rom[477][13] = 8'd24;
        rom[477][14] = -8'd14;
        rom[477][15] = 8'd30;
        rom[477][16] = 8'd31;
        rom[477][17] = 8'd4;
        rom[477][18] = -8'd9;
        rom[477][19] = -8'd11;
        rom[477][20] = -8'd6;
        rom[477][21] = 8'd37;
        rom[477][22] = -8'd38;
        rom[477][23] = 8'd24;
        rom[477][24] = -8'd3;
        rom[477][25] = 8'd9;
        rom[477][26] = -8'd12;
        rom[477][27] = -8'd46;
        rom[477][28] = -8'd7;
        rom[477][29] = 8'd16;
        rom[477][30] = -8'd21;
        rom[477][31] = 8'd39;
        rom[477][32] = 8'd10;
        rom[477][33] = 8'd24;
        rom[477][34] = 8'd12;
        rom[477][35] = -8'd1;
        rom[477][36] = 8'd0;
        rom[477][37] = -8'd50;
        rom[477][38] = -8'd53;
        rom[477][39] = -8'd18;
        rom[477][40] = -8'd13;
        rom[477][41] = -8'd4;
        rom[477][42] = 8'd2;
        rom[477][43] = -8'd4;
        rom[477][44] = -8'd16;
        rom[477][45] = 8'd2;
        rom[477][46] = 8'd19;
        rom[477][47] = -8'd50;
        rom[477][48] = -8'd74;
        rom[477][49] = -8'd10;
        rom[477][50] = 8'd12;
        rom[477][51] = -8'd1;
        rom[477][52] = 8'd24;
        rom[477][53] = 8'd40;
        rom[477][54] = 8'd0;
        rom[477][55] = 8'd19;
        rom[477][56] = -8'd21;
        rom[477][57] = 8'd3;
        rom[477][58] = -8'd6;
        rom[477][59] = -8'd1;
        rom[477][60] = -8'd8;
        rom[477][61] = 8'd8;
        rom[477][62] = 8'd3;
        rom[477][63] = -8'd3;
        rom[478][0] = 8'd9;
        rom[478][1] = -8'd20;
        rom[478][2] = 8'd32;
        rom[478][3] = 8'd12;
        rom[478][4] = 8'd18;
        rom[478][5] = 8'd11;
        rom[478][6] = 8'd20;
        rom[478][7] = -8'd35;
        rom[478][8] = -8'd4;
        rom[478][9] = -8'd15;
        rom[478][10] = 8'd7;
        rom[478][11] = 8'd14;
        rom[478][12] = 8'd11;
        rom[478][13] = -8'd16;
        rom[478][14] = -8'd45;
        rom[478][15] = -8'd19;
        rom[478][16] = -8'd39;
        rom[478][17] = -8'd32;
        rom[478][18] = -8'd25;
        rom[478][19] = 8'd10;
        rom[478][20] = -8'd11;
        rom[478][21] = 8'd14;
        rom[478][22] = -8'd5;
        rom[478][23] = 8'd27;
        rom[478][24] = -8'd10;
        rom[478][25] = 8'd15;
        rom[478][26] = -8'd33;
        rom[478][27] = 8'd13;
        rom[478][28] = 8'd11;
        rom[478][29] = -8'd8;
        rom[478][30] = -8'd1;
        rom[478][31] = -8'd33;
        rom[478][32] = 8'd6;
        rom[478][33] = 8'd2;
        rom[478][34] = -8'd4;
        rom[478][35] = 8'd13;
        rom[478][36] = -8'd47;
        rom[478][37] = 8'd1;
        rom[478][38] = -8'd20;
        rom[478][39] = 8'd2;
        rom[478][40] = 8'd16;
        rom[478][41] = 8'd5;
        rom[478][42] = -8'd12;
        rom[478][43] = 8'd2;
        rom[478][44] = 8'd30;
        rom[478][45] = -8'd33;
        rom[478][46] = -8'd12;
        rom[478][47] = -8'd28;
        rom[478][48] = -8'd4;
        rom[478][49] = -8'd4;
        rom[478][50] = 8'd32;
        rom[478][51] = -8'd36;
        rom[478][52] = 8'd25;
        rom[478][53] = -8'd4;
        rom[478][54] = -8'd20;
        rom[478][55] = 8'd1;
        rom[478][56] = -8'd34;
        rom[478][57] = -8'd30;
        rom[478][58] = 8'd16;
        rom[478][59] = -8'd3;
        rom[478][60] = 8'd29;
        rom[478][61] = -8'd7;
        rom[478][62] = 8'd9;
        rom[478][63] = -8'd3;
        rom[479][0] = 8'd11;
        rom[479][1] = -8'd9;
        rom[479][2] = -8'd34;
        rom[479][3] = 8'd8;
        rom[479][4] = -8'd33;
        rom[479][5] = 8'd13;
        rom[479][6] = -8'd87;
        rom[479][7] = -8'd2;
        rom[479][8] = -8'd23;
        rom[479][9] = 8'd19;
        rom[479][10] = 8'd37;
        rom[479][11] = -8'd12;
        rom[479][12] = 8'd0;
        rom[479][13] = 8'd25;
        rom[479][14] = 8'd16;
        rom[479][15] = 8'd26;
        rom[479][16] = 8'd4;
        rom[479][17] = 8'd2;
        rom[479][18] = -8'd1;
        rom[479][19] = -8'd7;
        rom[479][20] = -8'd6;
        rom[479][21] = 8'd38;
        rom[479][22] = -8'd14;
        rom[479][23] = 8'd23;
        rom[479][24] = 8'd23;
        rom[479][25] = -8'd3;
        rom[479][26] = 8'd48;
        rom[479][27] = 8'd2;
        rom[479][28] = 8'd15;
        rom[479][29] = 8'd11;
        rom[479][30] = 8'd22;
        rom[479][31] = 8'd6;
        rom[479][32] = -8'd7;
        rom[479][33] = -8'd25;
        rom[479][34] = 8'd12;
        rom[479][35] = -8'd5;
        rom[479][36] = 8'd0;
        rom[479][37] = 8'd3;
        rom[479][38] = 8'd11;
        rom[479][39] = -8'd2;
        rom[479][40] = 8'd31;
        rom[479][41] = 8'd2;
        rom[479][42] = -8'd16;
        rom[479][43] = -8'd7;
        rom[479][44] = -8'd13;
        rom[479][45] = -8'd55;
        rom[479][46] = -8'd37;
        rom[479][47] = -8'd15;
        rom[479][48] = 8'd6;
        rom[479][49] = 8'd11;
        rom[479][50] = 8'd7;
        rom[479][51] = -8'd35;
        rom[479][52] = 8'd31;
        rom[479][53] = -8'd2;
        rom[479][54] = 8'd8;
        rom[479][55] = -8'd31;
        rom[479][56] = 8'd36;
        rom[479][57] = 8'd0;
        rom[479][58] = 8'd24;
        rom[479][59] = 8'd9;
        rom[479][60] = -8'd21;
        rom[479][61] = -8'd1;
        rom[479][62] = 8'd26;
        rom[479][63] = 8'd13;
        rom[480][0] = 8'd3;
        rom[480][1] = 8'd30;
        rom[480][2] = -8'd28;
        rom[480][3] = -8'd15;
        rom[480][4] = -8'd3;
        rom[480][5] = 8'd19;
        rom[480][6] = 8'd33;
        rom[480][7] = 8'd7;
        rom[480][8] = -8'd21;
        rom[480][9] = 8'd12;
        rom[480][10] = 8'd6;
        rom[480][11] = 8'd12;
        rom[480][12] = 8'd2;
        rom[480][13] = -8'd46;
        rom[480][14] = 8'd0;
        rom[480][15] = -8'd37;
        rom[480][16] = -8'd32;
        rom[480][17] = -8'd1;
        rom[480][18] = -8'd10;
        rom[480][19] = 8'd20;
        rom[480][20] = 8'd0;
        rom[480][21] = 8'd4;
        rom[480][22] = -8'd28;
        rom[480][23] = 8'd10;
        rom[480][24] = 8'd25;
        rom[480][25] = -8'd41;
        rom[480][26] = 8'd36;
        rom[480][27] = -8'd14;
        rom[480][28] = -8'd24;
        rom[480][29] = -8'd20;
        rom[480][30] = 8'd2;
        rom[480][31] = 8'd11;
        rom[480][32] = -8'd42;
        rom[480][33] = -8'd32;
        rom[480][34] = 8'd16;
        rom[480][35] = 8'd12;
        rom[480][36] = 8'd8;
        rom[480][37] = -8'd8;
        rom[480][38] = -8'd24;
        rom[480][39] = -8'd2;
        rom[480][40] = -8'd14;
        rom[480][41] = -8'd2;
        rom[480][42] = -8'd15;
        rom[480][43] = 8'd4;
        rom[480][44] = -8'd24;
        rom[480][45] = 8'd27;
        rom[480][46] = -8'd96;
        rom[480][47] = -8'd16;
        rom[480][48] = -8'd4;
        rom[480][49] = -8'd3;
        rom[480][50] = -8'd15;
        rom[480][51] = 8'd1;
        rom[480][52] = -8'd28;
        rom[480][53] = -8'd12;
        rom[480][54] = 8'd19;
        rom[480][55] = -8'd16;
        rom[480][56] = -8'd16;
        rom[480][57] = -8'd2;
        rom[480][58] = 8'd14;
        rom[480][59] = -8'd16;
        rom[480][60] = -8'd2;
        rom[480][61] = -8'd5;
        rom[480][62] = -8'd6;
        rom[480][63] = -8'd17;
        rom[481][0] = -8'd1;
        rom[481][1] = -8'd41;
        rom[481][2] = -8'd3;
        rom[481][3] = -8'd22;
        rom[481][4] = -8'd103;
        rom[481][5] = -8'd12;
        rom[481][6] = -8'd14;
        rom[481][7] = 8'd0;
        rom[481][8] = -8'd31;
        rom[481][9] = -8'd53;
        rom[481][10] = 8'd23;
        rom[481][11] = 8'd22;
        rom[481][12] = -8'd20;
        rom[481][13] = 8'd3;
        rom[481][14] = -8'd51;
        rom[481][15] = 8'd8;
        rom[481][16] = 8'd61;
        rom[481][17] = -8'd17;
        rom[481][18] = 8'd20;
        rom[481][19] = 8'd48;
        rom[481][20] = -8'd4;
        rom[481][21] = -8'd21;
        rom[481][22] = -8'd38;
        rom[481][23] = -8'd6;
        rom[481][24] = -8'd13;
        rom[481][25] = -8'd17;
        rom[481][26] = -8'd30;
        rom[481][27] = 8'd25;
        rom[481][28] = 8'd21;
        rom[481][29] = 8'd14;
        rom[481][30] = -8'd12;
        rom[481][31] = -8'd7;
        rom[481][32] = 8'd51;
        rom[481][33] = 8'd43;
        rom[481][34] = -8'd28;
        rom[481][35] = -8'd61;
        rom[481][36] = -8'd12;
        rom[481][37] = -8'd32;
        rom[481][38] = -8'd38;
        rom[481][39] = -8'd24;
        rom[481][40] = 8'd27;
        rom[481][41] = 8'd20;
        rom[481][42] = 8'd10;
        rom[481][43] = 8'd22;
        rom[481][44] = -8'd38;
        rom[481][45] = -8'd28;
        rom[481][46] = 8'd20;
        rom[481][47] = 8'd44;
        rom[481][48] = -8'd36;
        rom[481][49] = -8'd8;
        rom[481][50] = 8'd20;
        rom[481][51] = -8'd27;
        rom[481][52] = 8'd1;
        rom[481][53] = -8'd3;
        rom[481][54] = -8'd49;
        rom[481][55] = 8'd7;
        rom[481][56] = 8'd45;
        rom[481][57] = 8'd2;
        rom[481][58] = -8'd1;
        rom[481][59] = 8'd18;
        rom[481][60] = 8'd5;
        rom[481][61] = 8'd7;
        rom[481][62] = 8'd15;
        rom[481][63] = 8'd6;
        rom[482][0] = 8'd3;
        rom[482][1] = -8'd26;
        rom[482][2] = -8'd73;
        rom[482][3] = -8'd20;
        rom[482][4] = -8'd11;
        rom[482][5] = -8'd18;
        rom[482][6] = -8'd19;
        rom[482][7] = 8'd24;
        rom[482][8] = -8'd12;
        rom[482][9] = -8'd21;
        rom[482][10] = 8'd8;
        rom[482][11] = -8'd3;
        rom[482][12] = 8'd10;
        rom[482][13] = 8'd19;
        rom[482][14] = 8'd20;
        rom[482][15] = -8'd5;
        rom[482][16] = -8'd26;
        rom[482][17] = 8'd3;
        rom[482][18] = -8'd12;
        rom[482][19] = 8'd17;
        rom[482][20] = -8'd7;
        rom[482][21] = 8'd12;
        rom[482][22] = 8'd27;
        rom[482][23] = 8'd9;
        rom[482][24] = 8'd24;
        rom[482][25] = -8'd20;
        rom[482][26] = 8'd13;
        rom[482][27] = 8'd25;
        rom[482][28] = -8'd16;
        rom[482][29] = 8'd22;
        rom[482][30] = 8'd7;
        rom[482][31] = -8'd50;
        rom[482][32] = -8'd51;
        rom[482][33] = 8'd37;
        rom[482][34] = 8'd2;
        rom[482][35] = 8'd11;
        rom[482][36] = 8'd2;
        rom[482][37] = -8'd35;
        rom[482][38] = -8'd17;
        rom[482][39] = 8'd7;
        rom[482][40] = -8'd46;
        rom[482][41] = 8'd2;
        rom[482][42] = 8'd4;
        rom[482][43] = -8'd10;
        rom[482][44] = -8'd21;
        rom[482][45] = 8'd10;
        rom[482][46] = 8'd0;
        rom[482][47] = 8'd24;
        rom[482][48] = -8'd8;
        rom[482][49] = -8'd6;
        rom[482][50] = 8'd2;
        rom[482][51] = 8'd29;
        rom[482][52] = 8'd24;
        rom[482][53] = 8'd28;
        rom[482][54] = 8'd15;
        rom[482][55] = -8'd21;
        rom[482][56] = 8'd9;
        rom[482][57] = 8'd4;
        rom[482][58] = -8'd32;
        rom[482][59] = 8'd5;
        rom[482][60] = -8'd22;
        rom[482][61] = 8'd46;
        rom[482][62] = 8'd6;
        rom[482][63] = -8'd4;
        rom[483][0] = -8'd53;
        rom[483][1] = -8'd9;
        rom[483][2] = -8'd35;
        rom[483][3] = -8'd18;
        rom[483][4] = -8'd2;
        rom[483][5] = -8'd35;
        rom[483][6] = -8'd6;
        rom[483][7] = 8'd4;
        rom[483][8] = 8'd20;
        rom[483][9] = -8'd15;
        rom[483][10] = -8'd83;
        rom[483][11] = -8'd2;
        rom[483][12] = 8'd4;
        rom[483][13] = -8'd11;
        rom[483][14] = 8'd8;
        rom[483][15] = 8'd7;
        rom[483][16] = -8'd17;
        rom[483][17] = -8'd7;
        rom[483][18] = -8'd47;
        rom[483][19] = 8'd3;
        rom[483][20] = -8'd9;
        rom[483][21] = -8'd51;
        rom[483][22] = -8'd12;
        rom[483][23] = 8'd26;
        rom[483][24] = -8'd15;
        rom[483][25] = -8'd36;
        rom[483][26] = -8'd41;
        rom[483][27] = 8'd7;
        rom[483][28] = 8'd16;
        rom[483][29] = -8'd27;
        rom[483][30] = -8'd19;
        rom[483][31] = 8'd13;
        rom[483][32] = 8'd16;
        rom[483][33] = 8'd21;
        rom[483][34] = -8'd22;
        rom[483][35] = -8'd19;
        rom[483][36] = 8'd16;
        rom[483][37] = -8'd39;
        rom[483][38] = -8'd29;
        rom[483][39] = -8'd19;
        rom[483][40] = -8'd36;
        rom[483][41] = 8'd40;
        rom[483][42] = -8'd11;
        rom[483][43] = -8'd7;
        rom[483][44] = 8'd4;
        rom[483][45] = -8'd38;
        rom[483][46] = -8'd56;
        rom[483][47] = 8'd12;
        rom[483][48] = 8'd0;
        rom[483][49] = -8'd21;
        rom[483][50] = -8'd36;
        rom[483][51] = -8'd15;
        rom[483][52] = 8'd18;
        rom[483][53] = -8'd8;
        rom[483][54] = 8'd2;
        rom[483][55] = -8'd6;
        rom[483][56] = -8'd5;
        rom[483][57] = 8'd1;
        rom[483][58] = -8'd34;
        rom[483][59] = -8'd40;
        rom[483][60] = -8'd5;
        rom[483][61] = 8'd2;
        rom[483][62] = 8'd26;
        rom[483][63] = -8'd37;
        rom[484][0] = -8'd18;
        rom[484][1] = -8'd66;
        rom[484][2] = 8'd10;
        rom[484][3] = -8'd18;
        rom[484][4] = -8'd69;
        rom[484][5] = -8'd1;
        rom[484][6] = 8'd16;
        rom[484][7] = -8'd38;
        rom[484][8] = -8'd22;
        rom[484][9] = -8'd40;
        rom[484][10] = 8'd12;
        rom[484][11] = 8'd8;
        rom[484][12] = -8'd51;
        rom[484][13] = -8'd35;
        rom[484][14] = -8'd23;
        rom[484][15] = -8'd10;
        rom[484][16] = -8'd6;
        rom[484][17] = -8'd16;
        rom[484][18] = 8'd7;
        rom[484][19] = -8'd48;
        rom[484][20] = -8'd1;
        rom[484][21] = 8'd2;
        rom[484][22] = -8'd19;
        rom[484][23] = -8'd50;
        rom[484][24] = 8'd4;
        rom[484][25] = 8'd5;
        rom[484][26] = 8'd15;
        rom[484][27] = -8'd37;
        rom[484][28] = 8'd2;
        rom[484][29] = 8'd6;
        rom[484][30] = 8'd28;
        rom[484][31] = -8'd68;
        rom[484][32] = -8'd22;
        rom[484][33] = 8'd3;
        rom[484][34] = 8'd11;
        rom[484][35] = -8'd26;
        rom[484][36] = 8'd15;
        rom[484][37] = -8'd13;
        rom[484][38] = -8'd41;
        rom[484][39] = -8'd6;
        rom[484][40] = 8'd35;
        rom[484][41] = -8'd26;
        rom[484][42] = -8'd19;
        rom[484][43] = -8'd41;
        rom[484][44] = -8'd17;
        rom[484][45] = -8'd38;
        rom[484][46] = -8'd58;
        rom[484][47] = 8'd8;
        rom[484][48] = -8'd8;
        rom[484][49] = 8'd31;
        rom[484][50] = 8'd1;
        rom[484][51] = 8'd7;
        rom[484][52] = -8'd49;
        rom[484][53] = -8'd21;
        rom[484][54] = -8'd11;
        rom[484][55] = -8'd9;
        rom[484][56] = -8'd11;
        rom[484][57] = -8'd11;
        rom[484][58] = 8'd14;
        rom[484][59] = -8'd42;
        rom[484][60] = -8'd26;
        rom[484][61] = -8'd16;
        rom[484][62] = 8'd7;
        rom[484][63] = 8'd23;
        rom[485][0] = 8'd20;
        rom[485][1] = -8'd41;
        rom[485][2] = -8'd104;
        rom[485][3] = 8'd7;
        rom[485][4] = -8'd9;
        rom[485][5] = -8'd22;
        rom[485][6] = 8'd21;
        rom[485][7] = 8'd9;
        rom[485][8] = -8'd4;
        rom[485][9] = -8'd1;
        rom[485][10] = 8'd10;
        rom[485][11] = 8'd33;
        rom[485][12] = -8'd12;
        rom[485][13] = -8'd6;
        rom[485][14] = -8'd15;
        rom[485][15] = -8'd9;
        rom[485][16] = 8'd4;
        rom[485][17] = -8'd41;
        rom[485][18] = 8'd3;
        rom[485][19] = -8'd70;
        rom[485][20] = -8'd1;
        rom[485][21] = -8'd26;
        rom[485][22] = -8'd3;
        rom[485][23] = 8'd1;
        rom[485][24] = -8'd36;
        rom[485][25] = 8'd30;
        rom[485][26] = 8'd31;
        rom[485][27] = -8'd91;
        rom[485][28] = 8'd11;
        rom[485][29] = 8'd8;
        rom[485][30] = -8'd59;
        rom[485][31] = 8'd19;
        rom[485][32] = 8'd7;
        rom[485][33] = -8'd15;
        rom[485][34] = 8'd11;
        rom[485][35] = -8'd22;
        rom[485][36] = 8'd7;
        rom[485][37] = -8'd14;
        rom[485][38] = -8'd14;
        rom[485][39] = -8'd40;
        rom[485][40] = -8'd16;
        rom[485][41] = 8'd24;
        rom[485][42] = -8'd30;
        rom[485][43] = -8'd46;
        rom[485][44] = -8'd3;
        rom[485][45] = -8'd10;
        rom[485][46] = -8'd52;
        rom[485][47] = 8'd20;
        rom[485][48] = 8'd15;
        rom[485][49] = 8'd32;
        rom[485][50] = -8'd12;
        rom[485][51] = -8'd18;
        rom[485][52] = 8'd34;
        rom[485][53] = 8'd35;
        rom[485][54] = -8'd17;
        rom[485][55] = -8'd16;
        rom[485][56] = -8'd74;
        rom[485][57] = 8'd7;
        rom[485][58] = 8'd11;
        rom[485][59] = -8'd15;
        rom[485][60] = 8'd9;
        rom[485][61] = 8'd35;
        rom[485][62] = 8'd21;
        rom[485][63] = -8'd26;
        rom[486][0] = -8'd37;
        rom[486][1] = -8'd29;
        rom[486][2] = -8'd24;
        rom[486][3] = 8'd14;
        rom[486][4] = 8'd15;
        rom[486][5] = -8'd38;
        rom[486][6] = -8'd54;
        rom[486][7] = 8'd8;
        rom[486][8] = -8'd40;
        rom[486][9] = -8'd61;
        rom[486][10] = -8'd15;
        rom[486][11] = -8'd5;
        rom[486][12] = 8'd34;
        rom[486][13] = 8'd10;
        rom[486][14] = -8'd27;
        rom[486][15] = 8'd2;
        rom[486][16] = 8'd11;
        rom[486][17] = -8'd21;
        rom[486][18] = -8'd26;
        rom[486][19] = -8'd22;
        rom[486][20] = 8'd3;
        rom[486][21] = -8'd28;
        rom[486][22] = -8'd1;
        rom[486][23] = 8'd27;
        rom[486][24] = -8'd31;
        rom[486][25] = -8'd26;
        rom[486][26] = -8'd7;
        rom[486][27] = -8'd37;
        rom[486][28] = 8'd5;
        rom[486][29] = -8'd11;
        rom[486][30] = -8'd3;
        rom[486][31] = -8'd1;
        rom[486][32] = 8'd8;
        rom[486][33] = -8'd16;
        rom[486][34] = -8'd13;
        rom[486][35] = -8'd6;
        rom[486][36] = -8'd6;
        rom[486][37] = -8'd46;
        rom[486][38] = -8'd20;
        rom[486][39] = -8'd21;
        rom[486][40] = 8'd39;
        rom[486][41] = 8'd49;
        rom[486][42] = -8'd3;
        rom[486][43] = 8'd19;
        rom[486][44] = -8'd25;
        rom[486][45] = 8'd22;
        rom[486][46] = 8'd16;
        rom[486][47] = -8'd25;
        rom[486][48] = -8'd28;
        rom[486][49] = -8'd25;
        rom[486][50] = 8'd29;
        rom[486][51] = 8'd22;
        rom[486][52] = -8'd1;
        rom[486][53] = -8'd35;
        rom[486][54] = -8'd30;
        rom[486][55] = -8'd46;
        rom[486][56] = 8'd9;
        rom[486][57] = 8'd7;
        rom[486][58] = 8'd45;
        rom[486][59] = -8'd7;
        rom[486][60] = -8'd13;
        rom[486][61] = 8'd14;
        rom[486][62] = -8'd43;
        rom[486][63] = 8'd0;
        rom[487][0] = -8'd18;
        rom[487][1] = 8'd3;
        rom[487][2] = -8'd27;
        rom[487][3] = 8'd44;
        rom[487][4] = -8'd6;
        rom[487][5] = -8'd1;
        rom[487][6] = 8'd20;
        rom[487][7] = -8'd12;
        rom[487][8] = -8'd9;
        rom[487][9] = -8'd13;
        rom[487][10] = -8'd20;
        rom[487][11] = 8'd16;
        rom[487][12] = 8'd15;
        rom[487][13] = -8'd27;
        rom[487][14] = -8'd12;
        rom[487][15] = -8'd23;
        rom[487][16] = -8'd33;
        rom[487][17] = -8'd27;
        rom[487][18] = 8'd19;
        rom[487][19] = -8'd19;
        rom[487][20] = -8'd12;
        rom[487][21] = -8'd26;
        rom[487][22] = 8'd3;
        rom[487][23] = -8'd20;
        rom[487][24] = 8'd1;
        rom[487][25] = -8'd27;
        rom[487][26] = 8'd5;
        rom[487][27] = -8'd1;
        rom[487][28] = -8'd14;
        rom[487][29] = -8'd38;
        rom[487][30] = 8'd9;
        rom[487][31] = 8'd4;
        rom[487][32] = -8'd58;
        rom[487][33] = 8'd4;
        rom[487][34] = 8'd10;
        rom[487][35] = 8'd19;
        rom[487][36] = -8'd1;
        rom[487][37] = 8'd30;
        rom[487][38] = -8'd4;
        rom[487][39] = 8'd9;
        rom[487][40] = -8'd8;
        rom[487][41] = 8'd10;
        rom[487][42] = 8'd20;
        rom[487][43] = 8'd5;
        rom[487][44] = 8'd7;
        rom[487][45] = 8'd22;
        rom[487][46] = -8'd11;
        rom[487][47] = -8'd32;
        rom[487][48] = -8'd37;
        rom[487][49] = -8'd1;
        rom[487][50] = 8'd23;
        rom[487][51] = -8'd17;
        rom[487][52] = 8'd23;
        rom[487][53] = 8'd10;
        rom[487][54] = 8'd14;
        rom[487][55] = -8'd21;
        rom[487][56] = 8'd18;
        rom[487][57] = 8'd26;
        rom[487][58] = -8'd15;
        rom[487][59] = -8'd28;
        rom[487][60] = 8'd2;
        rom[487][61] = -8'd4;
        rom[487][62] = 8'd15;
        rom[487][63] = -8'd22;
        rom[488][0] = -8'd8;
        rom[488][1] = 8'd92;
        rom[488][2] = -8'd3;
        rom[488][3] = 8'd7;
        rom[488][4] = 8'd7;
        rom[488][5] = 8'd5;
        rom[488][6] = 8'd2;
        rom[488][7] = -8'd27;
        rom[488][8] = 8'd5;
        rom[488][9] = 8'd35;
        rom[488][10] = -8'd69;
        rom[488][11] = 8'd19;
        rom[488][12] = -8'd23;
        rom[488][13] = 8'd1;
        rom[488][14] = 8'd26;
        rom[488][15] = -8'd18;
        rom[488][16] = -8'd30;
        rom[488][17] = 8'd2;
        rom[488][18] = 8'd18;
        rom[488][19] = -8'd5;
        rom[488][20] = -8'd1;
        rom[488][21] = -8'd27;
        rom[488][22] = 8'd9;
        rom[488][23] = -8'd40;
        rom[488][24] = -8'd13;
        rom[488][25] = -8'd23;
        rom[488][26] = -8'd8;
        rom[488][27] = -8'd64;
        rom[488][28] = -8'd24;
        rom[488][29] = -8'd3;
        rom[488][30] = 8'd35;
        rom[488][31] = -8'd25;
        rom[488][32] = 8'd10;
        rom[488][33] = -8'd32;
        rom[488][34] = -8'd29;
        rom[488][35] = 8'd3;
        rom[488][36] = 8'd45;
        rom[488][37] = -8'd27;
        rom[488][38] = 8'd54;
        rom[488][39] = -8'd12;
        rom[488][40] = -8'd2;
        rom[488][41] = -8'd27;
        rom[488][42] = 8'd4;
        rom[488][43] = 8'd0;
        rom[488][44] = 8'd19;
        rom[488][45] = 8'd39;
        rom[488][46] = -8'd33;
        rom[488][47] = -8'd4;
        rom[488][48] = 8'd19;
        rom[488][49] = -8'd9;
        rom[488][50] = -8'd72;
        rom[488][51] = 8'd27;
        rom[488][52] = -8'd5;
        rom[488][53] = 8'd5;
        rom[488][54] = 8'd5;
        rom[488][55] = 8'd18;
        rom[488][56] = 8'd37;
        rom[488][57] = -8'd11;
        rom[488][58] = 8'd24;
        rom[488][59] = -8'd43;
        rom[488][60] = 8'd15;
        rom[488][61] = 8'd2;
        rom[488][62] = 8'd3;
        rom[488][63] = 8'd8;
        rom[489][0] = -8'd65;
        rom[489][1] = 8'd33;
        rom[489][2] = 8'd5;
        rom[489][3] = -8'd8;
        rom[489][4] = -8'd96;
        rom[489][5] = -8'd30;
        rom[489][6] = 8'd38;
        rom[489][7] = -8'd110;
        rom[489][8] = 8'd27;
        rom[489][9] = 8'd12;
        rom[489][10] = -8'd46;
        rom[489][11] = -8'd65;
        rom[489][12] = 8'd1;
        rom[489][13] = -8'd24;
        rom[489][14] = 8'd18;
        rom[489][15] = -8'd48;
        rom[489][16] = -8'd33;
        rom[489][17] = -8'd21;
        rom[489][18] = 8'd3;
        rom[489][19] = -8'd35;
        rom[489][20] = -8'd4;
        rom[489][21] = -8'd16;
        rom[489][22] = 8'd9;
        rom[489][23] = -8'd67;
        rom[489][24] = -8'd2;
        rom[489][25] = 8'd55;
        rom[489][26] = 8'd23;
        rom[489][27] = -8'd13;
        rom[489][28] = 8'd6;
        rom[489][29] = 8'd20;
        rom[489][30] = -8'd43;
        rom[489][31] = 8'd52;
        rom[489][32] = 8'd11;
        rom[489][33] = -8'd11;
        rom[489][34] = 8'd4;
        rom[489][35] = -8'd32;
        rom[489][36] = 8'd58;
        rom[489][37] = -8'd38;
        rom[489][38] = -8'd19;
        rom[489][39] = 8'd0;
        rom[489][40] = -8'd60;
        rom[489][41] = 8'd50;
        rom[489][42] = -8'd3;
        rom[489][43] = -8'd2;
        rom[489][44] = 8'd13;
        rom[489][45] = -8'd100;
        rom[489][46] = -8'd4;
        rom[489][47] = -8'd50;
        rom[489][48] = -8'd21;
        rom[489][49] = 8'd38;
        rom[489][50] = 8'd31;
        rom[489][51] = -8'd2;
        rom[489][52] = 8'd11;
        rom[489][53] = 8'd23;
        rom[489][54] = -8'd17;
        rom[489][55] = 8'd20;
        rom[489][56] = -8'd25;
        rom[489][57] = 8'd46;
        rom[489][58] = -8'd12;
        rom[489][59] = 8'd2;
        rom[489][60] = 8'd15;
        rom[489][61] = -8'd20;
        rom[489][62] = -8'd24;
        rom[489][63] = -8'd24;
        rom[490][0] = 8'd30;
        rom[490][1] = -8'd43;
        rom[490][2] = -8'd9;
        rom[490][3] = 8'd40;
        rom[490][4] = 8'd6;
        rom[490][5] = -8'd22;
        rom[490][6] = 8'd11;
        rom[490][7] = 8'd9;
        rom[490][8] = -8'd9;
        rom[490][9] = -8'd2;
        rom[490][10] = -8'd27;
        rom[490][11] = 8'd25;
        rom[490][12] = -8'd6;
        rom[490][13] = -8'd18;
        rom[490][14] = 8'd7;
        rom[490][15] = -8'd6;
        rom[490][16] = -8'd3;
        rom[490][17] = -8'd56;
        rom[490][18] = 8'd22;
        rom[490][19] = 8'd15;
        rom[490][20] = 8'd5;
        rom[490][21] = 8'd26;
        rom[490][22] = 8'd12;
        rom[490][23] = 8'd22;
        rom[490][24] = -8'd3;
        rom[490][25] = -8'd31;
        rom[490][26] = 8'd7;
        rom[490][27] = -8'd21;
        rom[490][28] = 8'd11;
        rom[490][29] = -8'd3;
        rom[490][30] = -8'd5;
        rom[490][31] = 8'd34;
        rom[490][32] = 8'd28;
        rom[490][33] = 8'd43;
        rom[490][34] = 8'd2;
        rom[490][35] = -8'd13;
        rom[490][36] = 8'd15;
        rom[490][37] = -8'd20;
        rom[490][38] = -8'd11;
        rom[490][39] = -8'd3;
        rom[490][40] = -8'd2;
        rom[490][41] = 8'd26;
        rom[490][42] = -8'd10;
        rom[490][43] = -8'd24;
        rom[490][44] = 8'd8;
        rom[490][45] = -8'd53;
        rom[490][46] = 8'd3;
        rom[490][47] = -8'd45;
        rom[490][48] = 8'd26;
        rom[490][49] = 8'd8;
        rom[490][50] = 8'd15;
        rom[490][51] = 8'd38;
        rom[490][52] = -8'd15;
        rom[490][53] = 8'd27;
        rom[490][54] = -8'd19;
        rom[490][55] = -8'd7;
        rom[490][56] = -8'd31;
        rom[490][57] = 8'd6;
        rom[490][58] = -8'd11;
        rom[490][59] = -8'd9;
        rom[490][60] = 8'd16;
        rom[490][61] = -8'd29;
        rom[490][62] = -8'd9;
        rom[490][63] = -8'd9;
        rom[491][0] = -8'd22;
        rom[491][1] = -8'd6;
        rom[491][2] = 8'd4;
        rom[491][3] = -8'd50;
        rom[491][4] = -8'd38;
        rom[491][5] = 8'd1;
        rom[491][6] = 8'd9;
        rom[491][7] = -8'd3;
        rom[491][8] = 8'd0;
        rom[491][9] = 8'd11;
        rom[491][10] = 8'd33;
        rom[491][11] = 8'd33;
        rom[491][12] = -8'd7;
        rom[491][13] = -8'd19;
        rom[491][14] = -8'd11;
        rom[491][15] = 8'd1;
        rom[491][16] = 8'd30;
        rom[491][17] = -8'd25;
        rom[491][18] = -8'd4;
        rom[491][19] = -8'd2;
        rom[491][20] = -8'd12;
        rom[491][21] = -8'd19;
        rom[491][22] = -8'd9;
        rom[491][23] = -8'd40;
        rom[491][24] = -8'd34;
        rom[491][25] = 8'd11;
        rom[491][26] = 8'd15;
        rom[491][27] = 8'd10;
        rom[491][28] = 8'd6;
        rom[491][29] = -8'd22;
        rom[491][30] = 8'd7;
        rom[491][31] = 8'd10;
        rom[491][32] = -8'd33;
        rom[491][33] = -8'd6;
        rom[491][34] = -8'd7;
        rom[491][35] = 8'd1;
        rom[491][36] = -8'd14;
        rom[491][37] = -8'd16;
        rom[491][38] = 8'd54;
        rom[491][39] = 8'd13;
        rom[491][40] = -8'd5;
        rom[491][41] = -8'd15;
        rom[491][42] = 8'd26;
        rom[491][43] = 8'd6;
        rom[491][44] = 8'd23;
        rom[491][45] = 8'd22;
        rom[491][46] = 8'd23;
        rom[491][47] = 8'd6;
        rom[491][48] = -8'd41;
        rom[491][49] = 8'd19;
        rom[491][50] = 8'd32;
        rom[491][51] = -8'd10;
        rom[491][52] = -8'd22;
        rom[491][53] = -8'd27;
        rom[491][54] = -8'd7;
        rom[491][55] = 8'd12;
        rom[491][56] = 8'd15;
        rom[491][57] = -8'd70;
        rom[491][58] = -8'd34;
        rom[491][59] = 8'd22;
        rom[491][60] = -8'd22;
        rom[491][61] = 8'd26;
        rom[491][62] = -8'd7;
        rom[491][63] = 8'd33;
        rom[492][0] = -8'd12;
        rom[492][1] = 8'd8;
        rom[492][2] = -8'd58;
        rom[492][3] = 8'd46;
        rom[492][4] = -8'd4;
        rom[492][5] = -8'd5;
        rom[492][6] = -8'd3;
        rom[492][7] = 8'd12;
        rom[492][8] = -8'd25;
        rom[492][9] = -8'd24;
        rom[492][10] = 8'd32;
        rom[492][11] = 8'd9;
        rom[492][12] = -8'd36;
        rom[492][13] = -8'd60;
        rom[492][14] = -8'd26;
        rom[492][15] = -8'd13;
        rom[492][16] = -8'd4;
        rom[492][17] = -8'd21;
        rom[492][18] = 8'd18;
        rom[492][19] = -8'd57;
        rom[492][20] = 8'd5;
        rom[492][21] = 8'd10;
        rom[492][22] = 8'd0;
        rom[492][23] = -8'd10;
        rom[492][24] = -8'd15;
        rom[492][25] = -8'd37;
        rom[492][26] = -8'd5;
        rom[492][27] = -8'd30;
        rom[492][28] = -8'd15;
        rom[492][29] = -8'd6;
        rom[492][30] = 8'd6;
        rom[492][31] = 8'd5;
        rom[492][32] = -8'd28;
        rom[492][33] = -8'd6;
        rom[492][34] = 8'd12;
        rom[492][35] = -8'd13;
        rom[492][36] = 8'd16;
        rom[492][37] = 8'd16;
        rom[492][38] = 8'd21;
        rom[492][39] = 8'd12;
        rom[492][40] = 8'd38;
        rom[492][41] = -8'd34;
        rom[492][42] = -8'd3;
        rom[492][43] = 8'd4;
        rom[492][44] = 8'd8;
        rom[492][45] = 8'd23;
        rom[492][46] = -8'd48;
        rom[492][47] = -8'd5;
        rom[492][48] = -8'd37;
        rom[492][49] = 8'd20;
        rom[492][50] = 8'd11;
        rom[492][51] = -8'd5;
        rom[492][52] = -8'd8;
        rom[492][53] = 8'd33;
        rom[492][54] = 8'd14;
        rom[492][55] = 8'd18;
        rom[492][56] = -8'd53;
        rom[492][57] = -8'd13;
        rom[492][58] = 8'd2;
        rom[492][59] = 8'd12;
        rom[492][60] = 8'd14;
        rom[492][61] = 8'd9;
        rom[492][62] = 8'd42;
        rom[492][63] = 8'd4;
        rom[493][0] = 8'd21;
        rom[493][1] = -8'd13;
        rom[493][2] = -8'd44;
        rom[493][3] = 8'd8;
        rom[493][4] = 8'd40;
        rom[493][5] = -8'd35;
        rom[493][6] = -8'd35;
        rom[493][7] = -8'd3;
        rom[493][8] = -8'd36;
        rom[493][9] = 8'd4;
        rom[493][10] = -8'd2;
        rom[493][11] = -8'd9;
        rom[493][12] = -8'd12;
        rom[493][13] = -8'd2;
        rom[493][14] = -8'd25;
        rom[493][15] = -8'd7;
        rom[493][16] = -8'd49;
        rom[493][17] = 8'd19;
        rom[493][18] = 8'd25;
        rom[493][19] = -8'd97;
        rom[493][20] = 8'd1;
        rom[493][21] = -8'd32;
        rom[493][22] = 8'd11;
        rom[493][23] = -8'd77;
        rom[493][24] = 8'd22;
        rom[493][25] = -8'd25;
        rom[493][26] = -8'd44;
        rom[493][27] = 8'd15;
        rom[493][28] = -8'd11;
        rom[493][29] = -8'd35;
        rom[493][30] = -8'd21;
        rom[493][31] = -8'd44;
        rom[493][32] = -8'd16;
        rom[493][33] = -8'd31;
        rom[493][34] = 8'd42;
        rom[493][35] = 8'd5;
        rom[493][36] = -8'd4;
        rom[493][37] = -8'd2;
        rom[493][38] = -8'd10;
        rom[493][39] = 8'd8;
        rom[493][40] = -8'd41;
        rom[493][41] = -8'd3;
        rom[493][42] = -8'd10;
        rom[493][43] = -8'd37;
        rom[493][44] = 8'd1;
        rom[493][45] = -8'd8;
        rom[493][46] = -8'd56;
        rom[493][47] = 8'd40;
        rom[493][48] = 8'd13;
        rom[493][49] = 8'd3;
        rom[493][50] = -8'd47;
        rom[493][51] = 8'd8;
        rom[493][52] = 8'd27;
        rom[493][53] = -8'd30;
        rom[493][54] = -8'd38;
        rom[493][55] = 8'd33;
        rom[493][56] = -8'd8;
        rom[493][57] = -8'd30;
        rom[493][58] = -8'd49;
        rom[493][59] = -8'd19;
        rom[493][60] = -8'd1;
        rom[493][61] = 8'd16;
        rom[493][62] = -8'd6;
        rom[493][63] = -8'd1;
        rom[494][0] = -8'd23;
        rom[494][1] = -8'd42;
        rom[494][2] = 8'd12;
        rom[494][3] = -8'd27;
        rom[494][4] = 8'd23;
        rom[494][5] = -8'd25;
        rom[494][6] = 8'd20;
        rom[494][7] = -8'd29;
        rom[494][8] = 8'd9;
        rom[494][9] = 8'd9;
        rom[494][10] = -8'd91;
        rom[494][11] = -8'd22;
        rom[494][12] = -8'd7;
        rom[494][13] = -8'd26;
        rom[494][14] = -8'd33;
        rom[494][15] = -8'd7;
        rom[494][16] = -8'd117;
        rom[494][17] = -8'd21;
        rom[494][18] = -8'd20;
        rom[494][19] = 8'd29;
        rom[494][20] = -8'd3;
        rom[494][21] = -8'd18;
        rom[494][22] = -8'd17;
        rom[494][23] = -8'd1;
        rom[494][24] = 8'd23;
        rom[494][25] = -8'd66;
        rom[494][26] = 8'd12;
        rom[494][27] = -8'd13;
        rom[494][28] = 8'd25;
        rom[494][29] = 8'd17;
        rom[494][30] = -8'd1;
        rom[494][31] = -8'd61;
        rom[494][32] = 8'd55;
        rom[494][33] = -8'd48;
        rom[494][34] = -8'd22;
        rom[494][35] = 8'd21;
        rom[494][36] = 8'd13;
        rom[494][37] = -8'd20;
        rom[494][38] = 8'd20;
        rom[494][39] = -8'd8;
        rom[494][40] = -8'd30;
        rom[494][41] = 8'd2;
        rom[494][42] = -8'd10;
        rom[494][43] = -8'd11;
        rom[494][44] = -8'd28;
        rom[494][45] = -8'd45;
        rom[494][46] = -8'd32;
        rom[494][47] = -8'd27;
        rom[494][48] = -8'd35;
        rom[494][49] = -8'd1;
        rom[494][50] = -8'd27;
        rom[494][51] = 8'd11;
        rom[494][52] = 8'd0;
        rom[494][53] = 8'd11;
        rom[494][54] = 8'd18;
        rom[494][55] = 8'd35;
        rom[494][56] = 8'd3;
        rom[494][57] = 8'd2;
        rom[494][58] = 8'd0;
        rom[494][59] = -8'd54;
        rom[494][60] = -8'd5;
        rom[494][61] = -8'd13;
        rom[494][62] = -8'd11;
        rom[494][63] = -8'd11;
        rom[495][0] = -8'd31;
        rom[495][1] = 8'd60;
        rom[495][2] = -8'd59;
        rom[495][3] = 8'd10;
        rom[495][4] = 8'd22;
        rom[495][5] = 8'd1;
        rom[495][6] = 8'd10;
        rom[495][7] = 8'd43;
        rom[495][8] = -8'd24;
        rom[495][9] = -8'd12;
        rom[495][10] = 8'd32;
        rom[495][11] = -8'd39;
        rom[495][12] = -8'd12;
        rom[495][13] = 8'd24;
        rom[495][14] = 8'd32;
        rom[495][15] = -8'd47;
        rom[495][16] = -8'd58;
        rom[495][17] = -8'd1;
        rom[495][18] = -8'd25;
        rom[495][19] = 8'd2;
        rom[495][20] = -8'd2;
        rom[495][21] = 8'd33;
        rom[495][22] = -8'd2;
        rom[495][23] = 8'd30;
        rom[495][24] = 8'd31;
        rom[495][25] = -8'd9;
        rom[495][26] = -8'd27;
        rom[495][27] = 8'd11;
        rom[495][28] = -8'd16;
        rom[495][29] = -8'd18;
        rom[495][30] = 8'd18;
        rom[495][31] = 8'd14;
        rom[495][32] = -8'd4;
        rom[495][33] = 8'd7;
        rom[495][34] = 8'd96;
        rom[495][35] = 8'd40;
        rom[495][36] = 8'd22;
        rom[495][37] = 8'd44;
        rom[495][38] = 8'd26;
        rom[495][39] = 8'd20;
        rom[495][40] = -8'd63;
        rom[495][41] = -8'd25;
        rom[495][42] = -8'd21;
        rom[495][43] = 8'd1;
        rom[495][44] = -8'd6;
        rom[495][45] = 8'd31;
        rom[495][46] = -8'd31;
        rom[495][47] = 8'd2;
        rom[495][48] = 8'd21;
        rom[495][49] = 8'd45;
        rom[495][50] = 8'd10;
        rom[495][51] = -8'd1;
        rom[495][52] = -8'd29;
        rom[495][53] = 8'd7;
        rom[495][54] = -8'd12;
        rom[495][55] = -8'd20;
        rom[495][56] = 8'd18;
        rom[495][57] = 8'd38;
        rom[495][58] = 8'd19;
        rom[495][59] = -8'd55;
        rom[495][60] = 8'd32;
        rom[495][61] = -8'd6;
        rom[495][62] = -8'd5;
        rom[495][63] = 8'd10;
        rom[496][0] = 8'd0;
        rom[496][1] = -8'd8;
        rom[496][2] = -8'd72;
        rom[496][3] = -8'd4;
        rom[496][4] = -8'd30;
        rom[496][5] = -8'd11;
        rom[496][6] = 8'd38;
        rom[496][7] = 8'd9;
        rom[496][8] = 8'd9;
        rom[496][9] = -8'd44;
        rom[496][10] = -8'd11;
        rom[496][11] = -8'd23;
        rom[496][12] = 8'd31;
        rom[496][13] = 8'd13;
        rom[496][14] = 8'd29;
        rom[496][15] = 8'd12;
        rom[496][16] = -8'd8;
        rom[496][17] = 8'd21;
        rom[496][18] = 8'd15;
        rom[496][19] = -8'd3;
        rom[496][20] = -8'd11;
        rom[496][21] = 8'd25;
        rom[496][22] = 8'd57;
        rom[496][23] = -8'd54;
        rom[496][24] = 8'd28;
        rom[496][25] = 8'd31;
        rom[496][26] = -8'd10;
        rom[496][27] = 8'd20;
        rom[496][28] = -8'd23;
        rom[496][29] = 8'd6;
        rom[496][30] = 8'd9;
        rom[496][31] = -8'd16;
        rom[496][32] = 8'd54;
        rom[496][33] = -8'd11;
        rom[496][34] = -8'd10;
        rom[496][35] = -8'd17;
        rom[496][36] = 8'd4;
        rom[496][37] = -8'd39;
        rom[496][38] = 8'd46;
        rom[496][39] = 8'd0;
        rom[496][40] = 8'd30;
        rom[496][41] = -8'd7;
        rom[496][42] = -8'd64;
        rom[496][43] = 8'd1;
        rom[496][44] = -8'd32;
        rom[496][45] = -8'd48;
        rom[496][46] = 8'd12;
        rom[496][47] = 8'd4;
        rom[496][48] = 8'd8;
        rom[496][49] = -8'd2;
        rom[496][50] = -8'd29;
        rom[496][51] = -8'd58;
        rom[496][52] = -8'd65;
        rom[496][53] = 8'd2;
        rom[496][54] = -8'd37;
        rom[496][55] = 8'd6;
        rom[496][56] = -8'd27;
        rom[496][57] = -8'd12;
        rom[496][58] = 8'd37;
        rom[496][59] = -8'd25;
        rom[496][60] = -8'd14;
        rom[496][61] = -8'd5;
        rom[496][62] = 8'd16;
        rom[496][63] = -8'd12;
        rom[497][0] = -8'd8;
        rom[497][1] = -8'd2;
        rom[497][2] = -8'd3;
        rom[497][3] = 8'd7;
        rom[497][4] = 8'd21;
        rom[497][5] = -8'd24;
        rom[497][6] = -8'd21;
        rom[497][7] = 8'd0;
        rom[497][8] = 8'd1;
        rom[497][9] = -8'd21;
        rom[497][10] = 8'd24;
        rom[497][11] = 8'd32;
        rom[497][12] = 8'd16;
        rom[497][13] = 8'd48;
        rom[497][14] = -8'd10;
        rom[497][15] = -8'd45;
        rom[497][16] = -8'd19;
        rom[497][17] = 8'd6;
        rom[497][18] = 8'd18;
        rom[497][19] = 8'd27;
        rom[497][20] = -8'd3;
        rom[497][21] = -8'd18;
        rom[497][22] = -8'd24;
        rom[497][23] = 8'd16;
        rom[497][24] = 8'd26;
        rom[497][25] = -8'd23;
        rom[497][26] = 8'd19;
        rom[497][27] = -8'd3;
        rom[497][28] = -8'd4;
        rom[497][29] = -8'd5;
        rom[497][30] = -8'd24;
        rom[497][31] = -8'd18;
        rom[497][32] = 8'd16;
        rom[497][33] = -8'd26;
        rom[497][34] = 8'd2;
        rom[497][35] = 8'd14;
        rom[497][36] = 8'd33;
        rom[497][37] = 8'd2;
        rom[497][38] = -8'd5;
        rom[497][39] = -8'd19;
        rom[497][40] = 8'd23;
        rom[497][41] = -8'd5;
        rom[497][42] = -8'd24;
        rom[497][43] = -8'd9;
        rom[497][44] = 8'd27;
        rom[497][45] = 8'd15;
        rom[497][46] = -8'd16;
        rom[497][47] = 8'd15;
        rom[497][48] = -8'd26;
        rom[497][49] = 8'd4;
        rom[497][50] = -8'd44;
        rom[497][51] = -8'd36;
        rom[497][52] = -8'd30;
        rom[497][53] = -8'd7;
        rom[497][54] = -8'd24;
        rom[497][55] = -8'd23;
        rom[497][56] = 8'd17;
        rom[497][57] = 8'd19;
        rom[497][58] = 8'd13;
        rom[497][59] = 8'd14;
        rom[497][60] = 8'd3;
        rom[497][61] = -8'd4;
        rom[497][62] = -8'd12;
        rom[497][63] = 8'd10;
        rom[498][0] = -8'd3;
        rom[498][1] = 8'd5;
        rom[498][2] = 8'd39;
        rom[498][3] = 8'd8;
        rom[498][4] = 8'd10;
        rom[498][5] = 8'd7;
        rom[498][6] = -8'd24;
        rom[498][7] = 8'd21;
        rom[498][8] = -8'd4;
        rom[498][9] = 8'd29;
        rom[498][10] = -8'd36;
        rom[498][11] = 8'd7;
        rom[498][12] = 8'd14;
        rom[498][13] = 8'd42;
        rom[498][14] = -8'd55;
        rom[498][15] = 8'd30;
        rom[498][16] = -8'd14;
        rom[498][17] = -8'd6;
        rom[498][18] = 8'd20;
        rom[498][19] = 8'd7;
        rom[498][20] = -8'd5;
        rom[498][21] = -8'd22;
        rom[498][22] = 8'd7;
        rom[498][23] = 8'd4;
        rom[498][24] = -8'd13;
        rom[498][25] = -8'd27;
        rom[498][26] = -8'd69;
        rom[498][27] = 8'd27;
        rom[498][28] = 8'd17;
        rom[498][29] = -8'd17;
        rom[498][30] = -8'd27;
        rom[498][31] = -8'd1;
        rom[498][32] = 8'd10;
        rom[498][33] = -8'd15;
        rom[498][34] = 8'd32;
        rom[498][35] = -8'd3;
        rom[498][36] = -8'd12;
        rom[498][37] = -8'd48;
        rom[498][38] = -8'd8;
        rom[498][39] = -8'd15;
        rom[498][40] = 8'd9;
        rom[498][41] = 8'd5;
        rom[498][42] = -8'd28;
        rom[498][43] = 8'd12;
        rom[498][44] = 8'd6;
        rom[498][45] = -8'd78;
        rom[498][46] = 8'd35;
        rom[498][47] = 8'd29;
        rom[498][48] = -8'd2;
        rom[498][49] = 8'd22;
        rom[498][50] = 8'd10;
        rom[498][51] = -8'd30;
        rom[498][52] = -8'd5;
        rom[498][53] = -8'd9;
        rom[498][54] = 8'd22;
        rom[498][55] = 8'd5;
        rom[498][56] = 8'd2;
        rom[498][57] = -8'd13;
        rom[498][58] = -8'd22;
        rom[498][59] = -8'd49;
        rom[498][60] = 8'd1;
        rom[498][61] = 8'd3;
        rom[498][62] = 8'd10;
        rom[498][63] = 8'd19;
        rom[499][0] = 8'd1;
        rom[499][1] = -8'd12;
        rom[499][2] = 8'd9;
        rom[499][3] = 8'd9;
        rom[499][4] = -8'd67;
        rom[499][5] = -8'd36;
        rom[499][6] = -8'd41;
        rom[499][7] = 8'd3;
        rom[499][8] = -8'd2;
        rom[499][9] = -8'd8;
        rom[499][10] = 8'd31;
        rom[499][11] = 8'd4;
        rom[499][12] = 8'd7;
        rom[499][13] = 8'd11;
        rom[499][14] = -8'd18;
        rom[499][15] = -8'd30;
        rom[499][16] = -8'd5;
        rom[499][17] = 8'd12;
        rom[499][18] = 8'd9;
        rom[499][19] = 8'd13;
        rom[499][20] = 8'd2;
        rom[499][21] = 8'd33;
        rom[499][22] = -8'd20;
        rom[499][23] = -8'd25;
        rom[499][24] = 8'd1;
        rom[499][25] = 8'd8;
        rom[499][26] = -8'd8;
        rom[499][27] = 8'd50;
        rom[499][28] = 8'd3;
        rom[499][29] = -8'd32;
        rom[499][30] = -8'd43;
        rom[499][31] = -8'd34;
        rom[499][32] = -8'd30;
        rom[499][33] = -8'd18;
        rom[499][34] = -8'd13;
        rom[499][35] = -8'd28;
        rom[499][36] = -8'd2;
        rom[499][37] = -8'd50;
        rom[499][38] = -8'd28;
        rom[499][39] = -8'd1;
        rom[499][40] = -8'd15;
        rom[499][41] = -8'd10;
        rom[499][42] = -8'd65;
        rom[499][43] = 8'd12;
        rom[499][44] = -8'd20;
        rom[499][45] = 8'd22;
        rom[499][46] = -8'd26;
        rom[499][47] = 8'd53;
        rom[499][48] = 8'd20;
        rom[499][49] = -8'd16;
        rom[499][50] = -8'd2;
        rom[499][51] = 8'd15;
        rom[499][52] = -8'd1;
        rom[499][53] = -8'd19;
        rom[499][54] = -8'd15;
        rom[499][55] = -8'd5;
        rom[499][56] = -8'd45;
        rom[499][57] = -8'd50;
        rom[499][58] = 8'd9;
        rom[499][59] = 8'd15;
        rom[499][60] = 8'd1;
        rom[499][61] = -8'd11;
        rom[499][62] = 8'd2;
        rom[499][63] = 8'd1;
        rom[500][0] = -8'd1;
        rom[500][1] = -8'd7;
        rom[500][2] = -8'd10;
        rom[500][3] = -8'd54;
        rom[500][4] = 8'd4;
        rom[500][5] = 8'd2;
        rom[500][6] = 8'd16;
        rom[500][7] = 8'd17;
        rom[500][8] = -8'd12;
        rom[500][9] = 8'd7;
        rom[500][10] = 8'd29;
        rom[500][11] = 8'd14;
        rom[500][12] = -8'd35;
        rom[500][13] = 8'd40;
        rom[500][14] = -8'd15;
        rom[500][15] = -8'd15;
        rom[500][16] = 8'd3;
        rom[500][17] = 8'd10;
        rom[500][18] = -8'd6;
        rom[500][19] = -8'd27;
        rom[500][20] = -8'd2;
        rom[500][21] = 8'd34;
        rom[500][22] = -8'd75;
        rom[500][23] = 8'd8;
        rom[500][24] = -8'd28;
        rom[500][25] = -8'd18;
        rom[500][26] = 8'd0;
        rom[500][27] = 8'd36;
        rom[500][28] = 8'd20;
        rom[500][29] = 8'd14;
        rom[500][30] = 8'd16;
        rom[500][31] = 8'd1;
        rom[500][32] = 8'd2;
        rom[500][33] = 8'd22;
        rom[500][34] = -8'd8;
        rom[500][35] = -8'd23;
        rom[500][36] = 8'd9;
        rom[500][37] = 8'd64;
        rom[500][38] = -8'd27;
        rom[500][39] = 8'd26;
        rom[500][40] = 8'd20;
        rom[500][41] = -8'd36;
        rom[500][42] = -8'd24;
        rom[500][43] = -8'd12;
        rom[500][44] = 8'd12;
        rom[500][45] = 8'd6;
        rom[500][46] = 8'd16;
        rom[500][47] = -8'd2;
        rom[500][48] = -8'd25;
        rom[500][49] = 8'd6;
        rom[500][50] = 8'd10;
        rom[500][51] = 8'd5;
        rom[500][52] = 8'd25;
        rom[500][53] = -8'd12;
        rom[500][54] = 8'd4;
        rom[500][55] = 8'd7;
        rom[500][56] = 8'd25;
        rom[500][57] = -8'd37;
        rom[500][58] = 8'd21;
        rom[500][59] = -8'd28;
        rom[500][60] = -8'd62;
        rom[500][61] = -8'd3;
        rom[500][62] = 8'd32;
        rom[500][63] = -8'd34;
        rom[501][0] = 8'd33;
        rom[501][1] = -8'd29;
        rom[501][2] = 8'd9;
        rom[501][3] = -8'd15;
        rom[501][4] = 8'd28;
        rom[501][5] = 8'd5;
        rom[501][6] = 8'd4;
        rom[501][7] = 8'd17;
        rom[501][8] = 8'd4;
        rom[501][9] = -8'd20;
        rom[501][10] = -8'd42;
        rom[501][11] = -8'd29;
        rom[501][12] = -8'd43;
        rom[501][13] = 8'd27;
        rom[501][14] = 8'd4;
        rom[501][15] = -8'd14;
        rom[501][16] = 8'd24;
        rom[501][17] = -8'd55;
        rom[501][18] = -8'd2;
        rom[501][19] = -8'd34;
        rom[501][20] = -8'd5;
        rom[501][21] = 8'd12;
        rom[501][22] = 8'd32;
        rom[501][23] = 8'd2;
        rom[501][24] = 8'd20;
        rom[501][25] = 8'd28;
        rom[501][26] = 8'd3;
        rom[501][27] = -8'd16;
        rom[501][28] = -8'd32;
        rom[501][29] = -8'd15;
        rom[501][30] = 8'd8;
        rom[501][31] = -8'd2;
        rom[501][32] = 8'd2;
        rom[501][33] = 8'd5;
        rom[501][34] = -8'd4;
        rom[501][35] = -8'd17;
        rom[501][36] = -8'd14;
        rom[501][37] = 8'd4;
        rom[501][38] = -8'd23;
        rom[501][39] = -8'd20;
        rom[501][40] = 8'd29;
        rom[501][41] = -8'd19;
        rom[501][42] = 8'd31;
        rom[501][43] = 8'd35;
        rom[501][44] = -8'd4;
        rom[501][45] = -8'd39;
        rom[501][46] = 8'd36;
        rom[501][47] = -8'd42;
        rom[501][48] = 8'd28;
        rom[501][49] = -8'd18;
        rom[501][50] = 8'd4;
        rom[501][51] = 8'd22;
        rom[501][52] = 8'd3;
        rom[501][53] = 8'd44;
        rom[501][54] = 8'd17;
        rom[501][55] = -8'd29;
        rom[501][56] = -8'd42;
        rom[501][57] = -8'd44;
        rom[501][58] = -8'd22;
        rom[501][59] = 8'd19;
        rom[501][60] = 8'd12;
        rom[501][61] = 8'd17;
        rom[501][62] = -8'd3;
        rom[501][63] = -8'd24;
        rom[502][0] = -8'd5;
        rom[502][1] = 8'd8;
        rom[502][2] = -8'd5;
        rom[502][3] = 8'd8;
        rom[502][4] = 8'd2;
        rom[502][5] = 8'd8;
        rom[502][6] = -8'd6;
        rom[502][7] = -8'd8;
        rom[502][8] = 8'd2;
        rom[502][9] = 8'd10;
        rom[502][10] = 8'd0;
        rom[502][11] = -8'd10;
        rom[502][12] = -8'd1;
        rom[502][13] = 8'd5;
        rom[502][14] = 8'd6;
        rom[502][15] = -8'd2;
        rom[502][16] = -8'd2;
        rom[502][17] = 8'd1;
        rom[502][18] = 8'd2;
        rom[502][19] = 8'd4;
        rom[502][20] = 8'd2;
        rom[502][21] = 8'd1;
        rom[502][22] = 8'd3;
        rom[502][23] = -8'd9;
        rom[502][24] = 8'd6;
        rom[502][25] = 8'd4;
        rom[502][26] = -8'd4;
        rom[502][27] = 8'd5;
        rom[502][28] = 8'd1;
        rom[502][29] = -8'd7;
        rom[502][30] = -8'd4;
        rom[502][31] = 8'd7;
        rom[502][32] = -8'd8;
        rom[502][33] = 8'd8;
        rom[502][34] = -8'd1;
        rom[502][35] = -8'd16;
        rom[502][36] = -8'd1;
        rom[502][37] = 8'd7;
        rom[502][38] = 8'd5;
        rom[502][39] = -8'd4;
        rom[502][40] = 8'd4;
        rom[502][41] = 8'd6;
        rom[502][42] = 8'd6;
        rom[502][43] = -8'd9;
        rom[502][44] = -8'd3;
        rom[502][45] = -8'd11;
        rom[502][46] = -8'd1;
        rom[502][47] = -8'd4;
        rom[502][48] = 8'd3;
        rom[502][49] = -8'd7;
        rom[502][50] = 8'd6;
        rom[502][51] = 8'd10;
        rom[502][52] = -8'd3;
        rom[502][53] = 8'd2;
        rom[502][54] = -8'd6;
        rom[502][55] = -8'd11;
        rom[502][56] = -8'd8;
        rom[502][57] = -8'd7;
        rom[502][58] = 8'd14;
        rom[502][59] = 8'd7;
        rom[502][60] = 8'd10;
        rom[502][61] = 8'd4;
        rom[502][62] = 8'd14;
        rom[502][63] = 8'd7;
        rom[503][0] = -8'd51;
        rom[503][1] = -8'd21;
        rom[503][2] = -8'd96;
        rom[503][3] = -8'd31;
        rom[503][4] = -8'd62;
        rom[503][5] = -8'd2;
        rom[503][6] = -8'd17;
        rom[503][7] = 8'd12;
        rom[503][8] = -8'd44;
        rom[503][9] = 8'd4;
        rom[503][10] = -8'd28;
        rom[503][11] = -8'd27;
        rom[503][12] = -8'd6;
        rom[503][13] = 8'd17;
        rom[503][14] = -8'd52;
        rom[503][15] = -8'd44;
        rom[503][16] = 8'd3;
        rom[503][17] = -8'd24;
        rom[503][18] = -8'd38;
        rom[503][19] = -8'd48;
        rom[503][20] = -8'd16;
        rom[503][21] = 8'd5;
        rom[503][22] = -8'd81;
        rom[503][23] = 8'd16;
        rom[503][24] = -8'd16;
        rom[503][25] = -8'd3;
        rom[503][26] = -8'd1;
        rom[503][27] = -8'd47;
        rom[503][28] = -8'd43;
        rom[503][29] = -8'd17;
        rom[503][30] = -8'd2;
        rom[503][31] = -8'd11;
        rom[503][32] = -8'd40;
        rom[503][33] = -8'd10;
        rom[503][34] = 8'd24;
        rom[503][35] = 8'd5;
        rom[503][36] = -8'd9;
        rom[503][37] = -8'd7;
        rom[503][38] = -8'd36;
        rom[503][39] = 8'd11;
        rom[503][40] = 8'd36;
        rom[503][41] = -8'd20;
        rom[503][42] = -8'd35;
        rom[503][43] = 8'd3;
        rom[503][44] = 8'd12;
        rom[503][45] = 8'd5;
        rom[503][46] = -8'd60;
        rom[503][47] = -8'd4;
        rom[503][48] = -8'd22;
        rom[503][49] = -8'd18;
        rom[503][50] = -8'd33;
        rom[503][51] = -8'd2;
        rom[503][52] = -8'd13;
        rom[503][53] = 8'd7;
        rom[503][54] = -8'd39;
        rom[503][55] = -8'd44;
        rom[503][56] = -8'd6;
        rom[503][57] = 8'd29;
        rom[503][58] = 8'd3;
        rom[503][59] = -8'd4;
        rom[503][60] = -8'd48;
        rom[503][61] = 8'd9;
        rom[503][62] = 8'd30;
        rom[503][63] = -8'd5;
        rom[504][0] = -8'd36;
        rom[504][1] = -8'd47;
        rom[504][2] = -8'd3;
        rom[504][3] = 8'd5;
        rom[504][4] = -8'd62;
        rom[504][5] = -8'd23;
        rom[504][6] = -8'd3;
        rom[504][7] = -8'd18;
        rom[504][8] = -8'd20;
        rom[504][9] = -8'd38;
        rom[504][10] = 8'd11;
        rom[504][11] = -8'd17;
        rom[504][12] = 8'd2;
        rom[504][13] = -8'd10;
        rom[504][14] = -8'd62;
        rom[504][15] = -8'd44;
        rom[504][16] = -8'd4;
        rom[504][17] = -8'd10;
        rom[504][18] = -8'd46;
        rom[504][19] = 8'd22;
        rom[504][20] = -8'd11;
        rom[504][21] = 8'd34;
        rom[504][22] = -8'd37;
        rom[504][23] = 8'd29;
        rom[504][24] = 8'd29;
        rom[504][25] = -8'd60;
        rom[504][26] = -8'd11;
        rom[504][27] = -8'd32;
        rom[504][28] = 8'd7;
        rom[504][29] = -8'd5;
        rom[504][30] = 8'd25;
        rom[504][31] = -8'd92;
        rom[504][32] = 8'd13;
        rom[504][33] = -8'd33;
        rom[504][34] = -8'd20;
        rom[504][35] = -8'd14;
        rom[504][36] = -8'd20;
        rom[504][37] = 8'd0;
        rom[504][38] = 8'd31;
        rom[504][39] = -8'd1;
        rom[504][40] = 8'd30;
        rom[504][41] = 8'd11;
        rom[504][42] = -8'd17;
        rom[504][43] = -8'd19;
        rom[504][44] = -8'd7;
        rom[504][45] = -8'd8;
        rom[504][46] = -8'd33;
        rom[504][47] = 8'd27;
        rom[504][48] = 8'd5;
        rom[504][49] = -8'd3;
        rom[504][50] = -8'd30;
        rom[504][51] = -8'd23;
        rom[504][52] = -8'd14;
        rom[504][53] = -8'd11;
        rom[504][54] = 8'd3;
        rom[504][55] = -8'd12;
        rom[504][56] = -8'd35;
        rom[504][57] = -8'd12;
        rom[504][58] = 8'd9;
        rom[504][59] = 8'd25;
        rom[504][60] = -8'd39;
        rom[504][61] = 8'd3;
        rom[504][62] = 8'd14;
        rom[504][63] = 8'd4;
        rom[505][0] = -8'd5;
        rom[505][1] = 8'd45;
        rom[505][2] = 8'd28;
        rom[505][3] = 8'd2;
        rom[505][4] = 8'd23;
        rom[505][5] = 8'd6;
        rom[505][6] = -8'd9;
        rom[505][7] = 8'd0;
        rom[505][8] = -8'd25;
        rom[505][9] = 8'd9;
        rom[505][10] = -8'd7;
        rom[505][11] = 8'd20;
        rom[505][12] = 8'd36;
        rom[505][13] = -8'd4;
        rom[505][14] = -8'd5;
        rom[505][15] = -8'd3;
        rom[505][16] = -8'd12;
        rom[505][17] = 8'd29;
        rom[505][18] = 8'd8;
        rom[505][19] = -8'd38;
        rom[505][20] = -8'd10;
        rom[505][21] = -8'd37;
        rom[505][22] = -8'd68;
        rom[505][23] = 8'd44;
        rom[505][24] = 8'd17;
        rom[505][25] = -8'd36;
        rom[505][26] = 8'd5;
        rom[505][27] = 8'd19;
        rom[505][28] = -8'd11;
        rom[505][29] = -8'd32;
        rom[505][30] = 8'd38;
        rom[505][31] = -8'd3;
        rom[505][32] = -8'd31;
        rom[505][33] = -8'd11;
        rom[505][34] = 8'd48;
        rom[505][35] = 8'd19;
        rom[505][36] = -8'd20;
        rom[505][37] = 8'd15;
        rom[505][38] = -8'd14;
        rom[505][39] = 8'd4;
        rom[505][40] = -8'd22;
        rom[505][41] = 8'd0;
        rom[505][42] = 8'd22;
        rom[505][43] = -8'd11;
        rom[505][44] = 8'd10;
        rom[505][45] = -8'd49;
        rom[505][46] = -8'd9;
        rom[505][47] = -8'd70;
        rom[505][48] = -8'd42;
        rom[505][49] = 8'd23;
        rom[505][50] = -8'd11;
        rom[505][51] = -8'd62;
        rom[505][52] = 8'd20;
        rom[505][53] = -8'd35;
        rom[505][54] = 8'd2;
        rom[505][55] = -8'd27;
        rom[505][56] = 8'd8;
        rom[505][57] = -8'd40;
        rom[505][58] = 8'd18;
        rom[505][59] = 8'd4;
        rom[505][60] = -8'd2;
        rom[505][61] = 8'd12;
        rom[505][62] = 8'd18;
        rom[505][63] = -8'd1;
        rom[506][0] = 8'd19;
        rom[506][1] = 8'd37;
        rom[506][2] = 8'd29;
        rom[506][3] = -8'd7;
        rom[506][4] = 8'd1;
        rom[506][5] = 8'd10;
        rom[506][6] = -8'd19;
        rom[506][7] = -8'd45;
        rom[506][8] = 8'd16;
        rom[506][9] = -8'd45;
        rom[506][10] = 8'd71;
        rom[506][11] = -8'd37;
        rom[506][12] = -8'd12;
        rom[506][13] = -8'd8;
        rom[506][14] = 8'd11;
        rom[506][15] = -8'd6;
        rom[506][16] = 8'd15;
        rom[506][17] = 8'd21;
        rom[506][18] = 8'd39;
        rom[506][19] = -8'd19;
        rom[506][20] = -8'd7;
        rom[506][21] = -8'd17;
        rom[506][22] = -8'd6;
        rom[506][23] = 8'd3;
        rom[506][24] = -8'd19;
        rom[506][25] = 8'd27;
        rom[506][26] = -8'd6;
        rom[506][27] = -8'd4;
        rom[506][28] = 8'd11;
        rom[506][29] = -8'd27;
        rom[506][30] = 8'd16;
        rom[506][31] = 8'd23;
        rom[506][32] = 8'd5;
        rom[506][33] = 8'd20;
        rom[506][34] = 8'd0;
        rom[506][35] = -8'd82;
        rom[506][36] = 8'd15;
        rom[506][37] = 8'd33;
        rom[506][38] = -8'd61;
        rom[506][39] = -8'd9;
        rom[506][40] = -8'd32;
        rom[506][41] = 8'd25;
        rom[506][42] = 8'd27;
        rom[506][43] = 8'd3;
        rom[506][44] = -8'd10;
        rom[506][45] = -8'd13;
        rom[506][46] = 8'd13;
        rom[506][47] = -8'd13;
        rom[506][48] = 8'd15;
        rom[506][49] = 8'd26;
        rom[506][50] = -8'd74;
        rom[506][51] = 8'd28;
        rom[506][52] = -8'd31;
        rom[506][53] = 8'd35;
        rom[506][54] = 8'd30;
        rom[506][55] = 8'd14;
        rom[506][56] = 8'd37;
        rom[506][57] = -8'd4;
        rom[506][58] = 8'd5;
        rom[506][59] = 8'd18;
        rom[506][60] = 8'd7;
        rom[506][61] = 8'd10;
        rom[506][62] = -8'd29;
        rom[506][63] = 8'd3;
        rom[507][0] = -8'd3;
        rom[507][1] = 8'd3;
        rom[507][2] = -8'd47;
        rom[507][3] = -8'd47;
        rom[507][4] = -8'd78;
        rom[507][5] = -8'd22;
        rom[507][6] = -8'd23;
        rom[507][7] = -8'd2;
        rom[507][8] = 8'd13;
        rom[507][9] = 8'd12;
        rom[507][10] = 8'd9;
        rom[507][11] = 8'd10;
        rom[507][12] = -8'd1;
        rom[507][13] = 8'd46;
        rom[507][14] = -8'd3;
        rom[507][15] = 8'd3;
        rom[507][16] = 8'd29;
        rom[507][17] = 8'd10;
        rom[507][18] = -8'd17;
        rom[507][19] = -8'd20;
        rom[507][20] = -8'd8;
        rom[507][21] = -8'd40;
        rom[507][22] = 8'd5;
        rom[507][23] = 8'd5;
        rom[507][24] = 8'd13;
        rom[507][25] = -8'd25;
        rom[507][26] = -8'd11;
        rom[507][27] = 8'd7;
        rom[507][28] = -8'd48;
        rom[507][29] = -8'd21;
        rom[507][30] = 8'd18;
        rom[507][31] = -8'd14;
        rom[507][32] = 8'd15;
        rom[507][33] = 8'd14;
        rom[507][34] = -8'd47;
        rom[507][35] = -8'd6;
        rom[507][36] = -8'd34;
        rom[507][37] = 8'd17;
        rom[507][38] = -8'd2;
        rom[507][39] = -8'd27;
        rom[507][40] = 8'd18;
        rom[507][41] = -8'd53;
        rom[507][42] = 8'd23;
        rom[507][43] = -8'd36;
        rom[507][44] = -8'd10;
        rom[507][45] = 8'd13;
        rom[507][46] = -8'd3;
        rom[507][47] = -8'd10;
        rom[507][48] = 8'd7;
        rom[507][49] = 8'd38;
        rom[507][50] = 8'd1;
        rom[507][51] = 8'd10;
        rom[507][52] = -8'd23;
        rom[507][53] = -8'd52;
        rom[507][54] = -8'd16;
        rom[507][55] = -8'd61;
        rom[507][56] = 8'd12;
        rom[507][57] = -8'd21;
        rom[507][58] = 8'd0;
        rom[507][59] = -8'd23;
        rom[507][60] = -8'd9;
        rom[507][61] = -8'd2;
        rom[507][62] = 8'd24;
        rom[507][63] = -8'd10;
        rom[508][0] = 8'd27;
        rom[508][1] = 8'd39;
        rom[508][2] = -8'd9;
        rom[508][3] = -8'd17;
        rom[508][4] = -8'd21;
        rom[508][5] = -8'd43;
        rom[508][6] = -8'd3;
        rom[508][7] = 8'd10;
        rom[508][8] = 8'd27;
        rom[508][9] = -8'd36;
        rom[508][10] = -8'd13;
        rom[508][11] = 8'd15;
        rom[508][12] = -8'd54;
        rom[508][13] = -8'd49;
        rom[508][14] = -8'd51;
        rom[508][15] = 8'd21;
        rom[508][16] = 8'd39;
        rom[508][17] = -8'd9;
        rom[508][18] = 8'd5;
        rom[508][19] = 8'd13;
        rom[508][20] = 8'd1;
        rom[508][21] = -8'd14;
        rom[508][22] = -8'd14;
        rom[508][23] = -8'd48;
        rom[508][24] = 8'd38;
        rom[508][25] = 8'd19;
        rom[508][26] = -8'd16;
        rom[508][27] = -8'd44;
        rom[508][28] = -8'd34;
        rom[508][29] = -8'd10;
        rom[508][30] = -8'd11;
        rom[508][31] = -8'd9;
        rom[508][32] = 8'd27;
        rom[508][33] = 8'd5;
        rom[508][34] = -8'd64;
        rom[508][35] = -8'd7;
        rom[508][36] = 8'd26;
        rom[508][37] = 8'd10;
        rom[508][38] = 8'd43;
        rom[508][39] = 8'd32;
        rom[508][40] = 8'd46;
        rom[508][41] = 8'd21;
        rom[508][42] = -8'd5;
        rom[508][43] = 8'd27;
        rom[508][44] = -8'd4;
        rom[508][45] = 8'd24;
        rom[508][46] = -8'd21;
        rom[508][47] = 8'd13;
        rom[508][48] = -8'd46;
        rom[508][49] = -8'd38;
        rom[508][50] = -8'd27;
        rom[508][51] = 8'd6;
        rom[508][52] = -8'd38;
        rom[508][53] = -8'd79;
        rom[508][54] = -8'd9;
        rom[508][55] = 8'd13;
        rom[508][56] = 8'd8;
        rom[508][57] = -8'd27;
        rom[508][58] = 8'd18;
        rom[508][59] = -8'd32;
        rom[508][60] = -8'd11;
        rom[508][61] = -8'd8;
        rom[508][62] = 8'd6;
        rom[508][63] = 8'd23;
        rom[509][0] = 8'd4;
        rom[509][1] = 8'd8;
        rom[509][2] = 8'd2;
        rom[509][3] = -8'd42;
        rom[509][4] = 8'd26;
        rom[509][5] = -8'd6;
        rom[509][6] = -8'd80;
        rom[509][7] = -8'd3;
        rom[509][8] = -8'd72;
        rom[509][9] = -8'd3;
        rom[509][10] = 8'd3;
        rom[509][11] = -8'd7;
        rom[509][12] = 8'd16;
        rom[509][13] = 8'd14;
        rom[509][14] = -8'd37;
        rom[509][15] = -8'd26;
        rom[509][16] = -8'd18;
        rom[509][17] = -8'd34;
        rom[509][18] = 8'd44;
        rom[509][19] = 8'd2;
        rom[509][20] = 8'd2;
        rom[509][21] = -8'd23;
        rom[509][22] = -8'd34;
        rom[509][23] = 8'd35;
        rom[509][24] = 8'd7;
        rom[509][25] = -8'd8;
        rom[509][26] = 8'd1;
        rom[509][27] = -8'd1;
        rom[509][28] = 8'd19;
        rom[509][29] = 8'd15;
        rom[509][30] = -8'd7;
        rom[509][31] = -8'd34;
        rom[509][32] = -8'd6;
        rom[509][33] = -8'd23;
        rom[509][34] = 8'd24;
        rom[509][35] = 8'd5;
        rom[509][36] = 8'd7;
        rom[509][37] = -8'd32;
        rom[509][38] = -8'd39;
        rom[509][39] = 8'd9;
        rom[509][40] = 8'd6;
        rom[509][41] = 8'd9;
        rom[509][42] = 8'd35;
        rom[509][43] = 8'd8;
        rom[509][44] = 8'd34;
        rom[509][45] = -8'd37;
        rom[509][46] = 8'd6;
        rom[509][47] = -8'd16;
        rom[509][48] = -8'd23;
        rom[509][49] = 8'd43;
        rom[509][50] = 8'd0;
        rom[509][51] = -8'd8;
        rom[509][52] = -8'd3;
        rom[509][53] = 8'd2;
        rom[509][54] = -8'd11;
        rom[509][55] = 8'd5;
        rom[509][56] = -8'd6;
        rom[509][57] = -8'd33;
        rom[509][58] = -8'd25;
        rom[509][59] = 8'd17;
        rom[509][60] = -8'd9;
        rom[509][61] = -8'd4;
        rom[509][62] = -8'd44;
        rom[509][63] = 8'd9;
        rom[510][0] = 8'd33;
        rom[510][1] = -8'd37;
        rom[510][2] = 8'd8;
        rom[510][3] = -8'd17;
        rom[510][4] = -8'd32;
        rom[510][5] = 8'd7;
        rom[510][6] = -8'd66;
        rom[510][7] = -8'd17;
        rom[510][8] = -8'd41;
        rom[510][9] = -8'd51;
        rom[510][10] = -8'd4;
        rom[510][11] = 8'd28;
        rom[510][12] = -8'd16;
        rom[510][13] = 8'd18;
        rom[510][14] = -8'd15;
        rom[510][15] = 8'd24;
        rom[510][16] = 8'd13;
        rom[510][17] = 8'd53;
        rom[510][18] = -8'd6;
        rom[510][19] = 8'd21;
        rom[510][20] = -8'd5;
        rom[510][21] = 8'd23;
        rom[510][22] = 8'd4;
        rom[510][23] = 8'd15;
        rom[510][24] = -8'd6;
        rom[510][25] = -8'd55;
        rom[510][26] = 8'd20;
        rom[510][27] = -8'd8;
        rom[510][28] = -8'd56;
        rom[510][29] = -8'd7;
        rom[510][30] = -8'd28;
        rom[510][31] = -8'd30;
        rom[510][32] = -8'd4;
        rom[510][33] = 8'd27;
        rom[510][34] = -8'd15;
        rom[510][35] = -8'd26;
        rom[510][36] = 8'd25;
        rom[510][37] = -8'd36;
        rom[510][38] = -8'd35;
        rom[510][39] = 8'd38;
        rom[510][40] = -8'd17;
        rom[510][41] = -8'd38;
        rom[510][42] = 8'd38;
        rom[510][43] = -8'd51;
        rom[510][44] = -8'd40;
        rom[510][45] = -8'd10;
        rom[510][46] = 8'd19;
        rom[510][47] = -8'd61;
        rom[510][48] = -8'd34;
        rom[510][49] = -8'd57;
        rom[510][50] = 8'd11;
        rom[510][51] = -8'd56;
        rom[510][52] = -8'd2;
        rom[510][53] = -8'd25;
        rom[510][54] = -8'd85;
        rom[510][55] = 8'd0;
        rom[510][56] = -8'd8;
        rom[510][57] = -8'd18;
        rom[510][58] = -8'd7;
        rom[510][59] = -8'd13;
        rom[510][60] = -8'd46;
        rom[510][61] = -8'd49;
        rom[510][62] = -8'd26;
        rom[510][63] = -8'd7;
        rom[511][0] = 8'd23;
        rom[511][1] = 8'd38;
        rom[511][2] = -8'd2;
        rom[511][3] = 8'd17;
        rom[511][4] = 8'd10;
        rom[511][5] = 8'd18;
        rom[511][6] = 8'd24;
        rom[511][7] = -8'd89;
        rom[511][8] = 8'd37;
        rom[511][9] = 8'd11;
        rom[511][10] = -8'd49;
        rom[511][11] = 8'd37;
        rom[511][12] = -8'd38;
        rom[511][13] = -8'd38;
        rom[511][14] = -8'd7;
        rom[511][15] = 8'd17;
        rom[511][16] = -8'd88;
        rom[511][17] = -8'd2;
        rom[511][18] = 8'd29;
        rom[511][19] = -8'd16;
        rom[511][20] = -8'd6;
        rom[511][21] = -8'd14;
        rom[511][22] = 8'd20;
        rom[511][23] = -8'd12;
        rom[511][24] = -8'd37;
        rom[511][25] = -8'd13;
        rom[511][26] = 8'd21;
        rom[511][27] = 8'd13;
        rom[511][28] = 8'd3;
        rom[511][29] = 8'd18;
        rom[511][30] = -8'd33;
        rom[511][31] = 8'd10;
        rom[511][32] = 8'd15;
        rom[511][33] = 8'd31;
        rom[511][34] = -8'd7;
        rom[511][35] = 8'd30;
        rom[511][36] = 8'd11;
        rom[511][37] = -8'd11;
        rom[511][38] = -8'd22;
        rom[511][39] = 8'd9;
        rom[511][40] = 8'd15;
        rom[511][41] = 8'd21;
        rom[511][42] = -8'd7;
        rom[511][43] = -8'd15;
        rom[511][44] = 8'd25;
        rom[511][45] = -8'd14;
        rom[511][46] = -8'd26;
        rom[511][47] = -8'd45;
        rom[511][48] = -8'd2;
        rom[511][49] = -8'd8;
        rom[511][50] = 8'd10;
        rom[511][51] = -8'd10;
        rom[511][52] = 8'd27;
        rom[511][53] = 8'd53;
        rom[511][54] = -8'd54;
        rom[511][55] = 8'd38;
        rom[511][56] = 8'd8;
        rom[511][57] = -8'd26;
        rom[511][58] = -8'd3;
        rom[511][59] = -8'd55;
        rom[511][60] = -8'd3;
        rom[511][61] = -8'd15;
        rom[511][62] = 8'd24;
        rom[511][63] = -8'd28;
        rom[512][0] = 8'd11;
        rom[512][1] = -8'd27;
        rom[512][2] = -8'd10;
        rom[512][3] = -8'd33;
        rom[512][4] = -8'd25;
        rom[512][5] = -8'd28;
        rom[512][6] = 8'd19;
        rom[512][7] = 8'd21;
        rom[512][8] = -8'd7;
        rom[512][9] = 8'd41;
        rom[512][10] = -8'd53;
        rom[512][11] = 8'd9;
        rom[512][12] = 8'd4;
        rom[512][13] = 8'd6;
        rom[512][14] = -8'd26;
        rom[512][15] = 8'd24;
        rom[512][16] = 8'd4;
        rom[512][17] = 8'd18;
        rom[512][18] = 8'd13;
        rom[512][19] = 8'd34;
        rom[512][20] = 8'd3;
        rom[512][21] = 8'd31;
        rom[512][22] = 8'd2;
        rom[512][23] = -8'd39;
        rom[512][24] = -8'd1;
        rom[512][25] = 8'd30;
        rom[512][26] = -8'd35;
        rom[512][27] = -8'd37;
        rom[512][28] = 8'd11;
        rom[512][29] = 8'd11;
        rom[512][30] = 8'd10;
        rom[512][31] = -8'd8;
        rom[512][32] = -8'd34;
        rom[512][33] = 8'd32;
        rom[512][34] = 8'd53;
        rom[512][35] = -8'd33;
        rom[512][36] = -8'd26;
        rom[512][37] = -8'd27;
        rom[512][38] = -8'd28;
        rom[512][39] = 8'd22;
        rom[512][40] = -8'd21;
        rom[512][41] = 8'd0;
        rom[512][42] = 8'd24;
        rom[512][43] = -8'd9;
        rom[512][44] = 8'd2;
        rom[512][45] = 8'd3;
        rom[512][46] = 8'd9;
        rom[512][47] = 8'd16;
        rom[512][48] = -8'd16;
        rom[512][49] = -8'd3;
        rom[512][50] = 8'd10;
        rom[512][51] = -8'd3;
        rom[512][52] = 8'd25;
        rom[512][53] = 8'd23;
        rom[512][54] = 8'd41;
        rom[512][55] = 8'd44;
        rom[512][56] = 8'd4;
        rom[512][57] = 8'd3;
        rom[512][58] = -8'd24;
        rom[512][59] = 8'd10;
        rom[512][60] = 8'd26;
        rom[512][61] = -8'd20;
        rom[512][62] = -8'd26;
        rom[512][63] = 8'd5;
        rom[513][0] = 8'd38;
        rom[513][1] = -8'd9;
        rom[513][2] = -8'd63;
        rom[513][3] = -8'd56;
        rom[513][4] = 8'd11;
        rom[513][5] = 8'd22;
        rom[513][6] = 8'd44;
        rom[513][7] = 8'd14;
        rom[513][8] = -8'd32;
        rom[513][9] = -8'd29;
        rom[513][10] = -8'd14;
        rom[513][11] = -8'd4;
        rom[513][12] = 8'd34;
        rom[513][13] = -8'd67;
        rom[513][14] = -8'd17;
        rom[513][15] = -8'd2;
        rom[513][16] = -8'd7;
        rom[513][17] = -8'd96;
        rom[513][18] = 8'd11;
        rom[513][19] = -8'd50;
        rom[513][20] = 8'd2;
        rom[513][21] = -8'd44;
        rom[513][22] = -8'd48;
        rom[513][23] = 8'd7;
        rom[513][24] = -8'd45;
        rom[513][25] = 8'd19;
        rom[513][26] = 8'd26;
        rom[513][27] = -8'd32;
        rom[513][28] = -8'd8;
        rom[513][29] = 8'd25;
        rom[513][30] = 8'd15;
        rom[513][31] = -8'd16;
        rom[513][32] = 8'd41;
        rom[513][33] = 8'd12;
        rom[513][34] = -8'd34;
        rom[513][35] = -8'd12;
        rom[513][36] = -8'd8;
        rom[513][37] = 8'd5;
        rom[513][38] = 8'd1;
        rom[513][39] = 8'd18;
        rom[513][40] = -8'd11;
        rom[513][41] = -8'd8;
        rom[513][42] = -8'd17;
        rom[513][43] = 8'd5;
        rom[513][44] = 8'd10;
        rom[513][45] = -8'd36;
        rom[513][46] = -8'd42;
        rom[513][47] = 8'd5;
        rom[513][48] = -8'd52;
        rom[513][49] = -8'd32;
        rom[513][50] = 8'd19;
        rom[513][51] = -8'd42;
        rom[513][52] = -8'd52;
        rom[513][53] = -8'd6;
        rom[513][54] = -8'd25;
        rom[513][55] = 8'd36;
        rom[513][56] = -8'd35;
        rom[513][57] = 8'd0;
        rom[513][58] = 8'd62;
        rom[513][59] = -8'd3;
        rom[513][60] = 8'd28;
        rom[513][61] = 8'd3;
        rom[513][62] = 8'd33;
        rom[513][63] = -8'd16;
        rom[514][0] = -8'd55;
        rom[514][1] = -8'd19;
        rom[514][2] = -8'd15;
        rom[514][3] = -8'd9;
        rom[514][4] = -8'd58;
        rom[514][5] = 8'd39;
        rom[514][6] = -8'd33;
        rom[514][7] = 8'd11;
        rom[514][8] = -8'd7;
        rom[514][9] = -8'd2;
        rom[514][10] = -8'd20;
        rom[514][11] = 8'd16;
        rom[514][12] = -8'd13;
        rom[514][13] = -8'd53;
        rom[514][14] = 8'd31;
        rom[514][15] = -8'd57;
        rom[514][16] = 8'd4;
        rom[514][17] = -8'd9;
        rom[514][18] = -8'd4;
        rom[514][19] = -8'd32;
        rom[514][20] = -8'd3;
        rom[514][21] = 8'd44;
        rom[514][22] = -8'd113;
        rom[514][23] = -8'd16;
        rom[514][24] = -8'd2;
        rom[514][25] = -8'd25;
        rom[514][26] = 8'd0;
        rom[514][27] = -8'd5;
        rom[514][28] = 8'd15;
        rom[514][29] = -8'd2;
        rom[514][30] = 8'd1;
        rom[514][31] = 8'd2;
        rom[514][32] = -8'd84;
        rom[514][33] = -8'd27;
        rom[514][34] = -8'd14;
        rom[514][35] = -8'd22;
        rom[514][36] = 8'd51;
        rom[514][37] = -8'd10;
        rom[514][38] = -8'd3;
        rom[514][39] = 8'd0;
        rom[514][40] = 8'd27;
        rom[514][41] = -8'd42;
        rom[514][42] = -8'd24;
        rom[514][43] = 8'd21;
        rom[514][44] = 8'd15;
        rom[514][45] = 8'd8;
        rom[514][46] = -8'd37;
        rom[514][47] = 8'd30;
        rom[514][48] = -8'd57;
        rom[514][49] = -8'd41;
        rom[514][50] = 8'd45;
        rom[514][51] = -8'd74;
        rom[514][52] = 8'd2;
        rom[514][53] = -8'd72;
        rom[514][54] = -8'd99;
        rom[514][55] = 8'd41;
        rom[514][56] = -8'd52;
        rom[514][57] = -8'd12;
        rom[514][58] = 8'd15;
        rom[514][59] = -8'd1;
        rom[514][60] = -8'd18;
        rom[514][61] = 8'd29;
        rom[514][62] = 8'd35;
        rom[514][63] = -8'd20;
        rom[515][0] = -8'd8;
        rom[515][1] = 8'd33;
        rom[515][2] = -8'd74;
        rom[515][3] = -8'd20;
        rom[515][4] = 8'd1;
        rom[515][5] = -8'd2;
        rom[515][6] = 8'd10;
        rom[515][7] = 8'd41;
        rom[515][8] = -8'd4;
        rom[515][9] = 8'd18;
        rom[515][10] = -8'd83;
        rom[515][11] = -8'd5;
        rom[515][12] = -8'd58;
        rom[515][13] = -8'd57;
        rom[515][14] = 8'd67;
        rom[515][15] = 8'd24;
        rom[515][16] = -8'd52;
        rom[515][17] = 8'd8;
        rom[515][18] = 8'd9;
        rom[515][19] = 8'd6;
        rom[515][20] = -8'd11;
        rom[515][21] = 8'd27;
        rom[515][22] = 8'd33;
        rom[515][23] = -8'd12;
        rom[515][24] = 8'd6;
        rom[515][25] = 8'd2;
        rom[515][26] = 8'd24;
        rom[515][27] = -8'd7;
        rom[515][28] = -8'd14;
        rom[515][29] = 8'd26;
        rom[515][30] = 8'd41;
        rom[515][31] = -8'd13;
        rom[515][32] = 8'd14;
        rom[515][33] = -8'd3;
        rom[515][34] = -8'd3;
        rom[515][35] = 8'd11;
        rom[515][36] = 8'd11;
        rom[515][37] = -8'd35;
        rom[515][38] = -8'd12;
        rom[515][39] = 8'd12;
        rom[515][40] = 8'd4;
        rom[515][41] = 8'd18;
        rom[515][42] = -8'd26;
        rom[515][43] = 8'd23;
        rom[515][44] = -8'd30;
        rom[515][45] = 8'd9;
        rom[515][46] = -8'd57;
        rom[515][47] = -8'd68;
        rom[515][48] = 8'd16;
        rom[515][49] = -8'd16;
        rom[515][50] = 8'd6;
        rom[515][51] = 8'd25;
        rom[515][52] = -8'd2;
        rom[515][53] = -8'd11;
        rom[515][54] = 8'd1;
        rom[515][55] = -8'd28;
        rom[515][56] = -8'd9;
        rom[515][57] = -8'd43;
        rom[515][58] = 8'd15;
        rom[515][59] = -8'd5;
        rom[515][60] = 8'd17;
        rom[515][61] = 8'd21;
        rom[515][62] = -8'd2;
        rom[515][63] = 8'd2;
        rom[516][0] = -8'd70;
        rom[516][1] = -8'd47;
        rom[516][2] = -8'd46;
        rom[516][3] = 8'd16;
        rom[516][4] = 8'd39;
        rom[516][5] = -8'd34;
        rom[516][6] = -8'd79;
        rom[516][7] = -8'd36;
        rom[516][8] = 8'd5;
        rom[516][9] = -8'd16;
        rom[516][10] = -8'd56;
        rom[516][11] = 8'd8;
        rom[516][12] = -8'd15;
        rom[516][13] = -8'd20;
        rom[516][14] = -8'd32;
        rom[516][15] = -8'd6;
        rom[516][16] = 8'd34;
        rom[516][17] = 8'd1;
        rom[516][18] = 8'd14;
        rom[516][19] = 8'd1;
        rom[516][20] = 8'd0;
        rom[516][21] = -8'd66;
        rom[516][22] = -8'd26;
        rom[516][23] = -8'd22;
        rom[516][24] = -8'd20;
        rom[516][25] = -8'd1;
        rom[516][26] = -8'd29;
        rom[516][27] = -8'd43;
        rom[516][28] = -8'd15;
        rom[516][29] = -8'd12;
        rom[516][30] = 8'd19;
        rom[516][31] = -8'd24;
        rom[516][32] = 8'd39;
        rom[516][33] = -8'd8;
        rom[516][34] = 8'd0;
        rom[516][35] = -8'd59;
        rom[516][36] = -8'd23;
        rom[516][37] = 8'd23;
        rom[516][38] = -8'd15;
        rom[516][39] = -8'd28;
        rom[516][40] = -8'd28;
        rom[516][41] = 8'd39;
        rom[516][42] = 8'd27;
        rom[516][43] = -8'd22;
        rom[516][44] = 8'd4;
        rom[516][45] = -8'd3;
        rom[516][46] = -8'd29;
        rom[516][47] = -8'd26;
        rom[516][48] = -8'd60;
        rom[516][49] = -8'd66;
        rom[516][50] = -8'd14;
        rom[516][51] = 8'd3;
        rom[516][52] = -8'd68;
        rom[516][53] = -8'd32;
        rom[516][54] = -8'd8;
        rom[516][55] = -8'd41;
        rom[516][56] = -8'd5;
        rom[516][57] = 8'd14;
        rom[516][58] = -8'd15;
        rom[516][59] = -8'd32;
        rom[516][60] = 8'd19;
        rom[516][61] = -8'd15;
        rom[516][62] = -8'd20;
        rom[516][63] = -8'd15;
        rom[517][0] = 8'd8;
        rom[517][1] = -8'd1;
        rom[517][2] = -8'd2;
        rom[517][3] = -8'd6;
        rom[517][4] = 8'd4;
        rom[517][5] = -8'd3;
        rom[517][6] = -8'd2;
        rom[517][7] = -8'd8;
        rom[517][8] = -8'd4;
        rom[517][9] = -8'd2;
        rom[517][10] = 8'd7;
        rom[517][11] = 8'd5;
        rom[517][12] = -8'd6;
        rom[517][13] = 8'd2;
        rom[517][14] = -8'd3;
        rom[517][15] = 8'd0;
        rom[517][16] = -8'd8;
        rom[517][17] = -8'd3;
        rom[517][18] = 8'd7;
        rom[517][19] = 8'd7;
        rom[517][20] = 8'd9;
        rom[517][21] = -8'd4;
        rom[517][22] = -8'd8;
        rom[517][23] = 8'd8;
        rom[517][24] = -8'd7;
        rom[517][25] = 8'd1;
        rom[517][26] = 8'd10;
        rom[517][27] = -8'd6;
        rom[517][28] = 8'd0;
        rom[517][29] = -8'd3;
        rom[517][30] = -8'd11;
        rom[517][31] = 8'd1;
        rom[517][32] = 8'd7;
        rom[517][33] = 8'd1;
        rom[517][34] = -8'd9;
        rom[517][35] = 8'd2;
        rom[517][36] = -8'd5;
        rom[517][37] = 8'd5;
        rom[517][38] = 8'd1;
        rom[517][39] = 8'd2;
        rom[517][40] = 8'd4;
        rom[517][41] = 8'd7;
        rom[517][42] = 8'd8;
        rom[517][43] = -8'd1;
        rom[517][44] = 8'd1;
        rom[517][45] = 8'd4;
        rom[517][46] = -8'd1;
        rom[517][47] = 8'd7;
        rom[517][48] = -8'd6;
        rom[517][49] = 8'd2;
        rom[517][50] = 8'd1;
        rom[517][51] = -8'd5;
        rom[517][52] = -8'd2;
        rom[517][53] = -8'd2;
        rom[517][54] = -8'd4;
        rom[517][55] = 8'd1;
        rom[517][56] = -8'd4;
        rom[517][57] = 8'd1;
        rom[517][58] = 8'd1;
        rom[517][59] = 8'd2;
        rom[517][60] = 8'd8;
        rom[517][61] = 8'd1;
        rom[517][62] = 8'd7;
        rom[517][63] = 8'd10;
        rom[518][0] = -8'd16;
        rom[518][1] = -8'd22;
        rom[518][2] = -8'd4;
        rom[518][3] = 8'd38;
        rom[518][4] = -8'd37;
        rom[518][5] = -8'd7;
        rom[518][6] = -8'd28;
        rom[518][7] = 8'd21;
        rom[518][8] = 8'd45;
        rom[518][9] = 8'd10;
        rom[518][10] = -8'd43;
        rom[518][11] = 8'd23;
        rom[518][12] = -8'd87;
        rom[518][13] = -8'd7;
        rom[518][14] = -8'd31;
        rom[518][15] = -8'd3;
        rom[518][16] = -8'd30;
        rom[518][17] = 8'd68;
        rom[518][18] = 8'd35;
        rom[518][19] = -8'd22;
        rom[518][20] = 8'd0;
        rom[518][21] = 8'd13;
        rom[518][22] = -8'd33;
        rom[518][23] = 8'd31;
        rom[518][24] = -8'd8;
        rom[518][25] = -8'd36;
        rom[518][26] = -8'd15;
        rom[518][27] = 8'd25;
        rom[518][28] = 8'd28;
        rom[518][29] = -8'd10;
        rom[518][30] = 8'd44;
        rom[518][31] = 8'd15;
        rom[518][32] = -8'd29;
        rom[518][33] = -8'd9;
        rom[518][34] = 8'd43;
        rom[518][35] = 8'd23;
        rom[518][36] = -8'd65;
        rom[518][37] = -8'd32;
        rom[518][38] = -8'd16;
        rom[518][39] = -8'd17;
        rom[518][40] = 8'd7;
        rom[518][41] = -8'd14;
        rom[518][42] = 8'd19;
        rom[518][43] = -8'd43;
        rom[518][44] = -8'd46;
        rom[518][45] = -8'd18;
        rom[518][46] = -8'd14;
        rom[518][47] = 8'd35;
        rom[518][48] = 8'd43;
        rom[518][49] = -8'd24;
        rom[518][50] = -8'd5;
        rom[518][51] = -8'd10;
        rom[518][52] = -8'd21;
        rom[518][53] = -8'd1;
        rom[518][54] = 8'd31;
        rom[518][55] = -8'd74;
        rom[518][56] = 8'd5;
        rom[518][57] = -8'd11;
        rom[518][58] = 8'd5;
        rom[518][59] = 8'd12;
        rom[518][60] = -8'd23;
        rom[518][61] = -8'd26;
        rom[518][62] = 8'd21;
        rom[518][63] = 8'd1;
        rom[519][0] = 8'd27;
        rom[519][1] = 8'd18;
        rom[519][2] = -8'd17;
        rom[519][3] = 8'd26;
        rom[519][4] = 8'd6;
        rom[519][5] = 8'd15;
        rom[519][6] = -8'd30;
        rom[519][7] = -8'd14;
        rom[519][8] = 8'd16;
        rom[519][9] = -8'd22;
        rom[519][10] = -8'd17;
        rom[519][11] = -8'd24;
        rom[519][12] = 8'd18;
        rom[519][13] = 8'd23;
        rom[519][14] = -8'd12;
        rom[519][15] = 8'd23;
        rom[519][16] = -8'd2;
        rom[519][17] = -8'd10;
        rom[519][18] = 8'd34;
        rom[519][19] = -8'd22;
        rom[519][20] = 8'd2;
        rom[519][21] = 8'd2;
        rom[519][22] = 8'd25;
        rom[519][23] = 8'd25;
        rom[519][24] = -8'd40;
        rom[519][25] = 8'd15;
        rom[519][26] = 8'd13;
        rom[519][27] = 8'd17;
        rom[519][28] = 8'd23;
        rom[519][29] = -8'd3;
        rom[519][30] = -8'd44;
        rom[519][31] = -8'd42;
        rom[519][32] = 8'd20;
        rom[519][33] = -8'd42;
        rom[519][34] = 8'd6;
        rom[519][35] = 8'd16;
        rom[519][36] = 8'd21;
        rom[519][37] = -8'd31;
        rom[519][38] = -8'd30;
        rom[519][39] = -8'd35;
        rom[519][40] = 8'd25;
        rom[519][41] = -8'd13;
        rom[519][42] = 8'd6;
        rom[519][43] = 8'd1;
        rom[519][44] = 8'd7;
        rom[519][45] = -8'd23;
        rom[519][46] = -8'd13;
        rom[519][47] = -8'd27;
        rom[519][48] = 8'd10;
        rom[519][49] = -8'd31;
        rom[519][50] = -8'd22;
        rom[519][51] = -8'd71;
        rom[519][52] = -8'd69;
        rom[519][53] = -8'd26;
        rom[519][54] = 8'd5;
        rom[519][55] = -8'd15;
        rom[519][56] = -8'd22;
        rom[519][57] = 8'd31;
        rom[519][58] = -8'd18;
        rom[519][59] = -8'd27;
        rom[519][60] = -8'd27;
        rom[519][61] = -8'd49;
        rom[519][62] = 8'd9;
        rom[519][63] = 8'd14;
        rom[520][0] = 8'd1;
        rom[520][1] = -8'd1;
        rom[520][2] = 8'd32;
        rom[520][3] = -8'd5;
        rom[520][4] = 8'd10;
        rom[520][5] = 8'd1;
        rom[520][6] = -8'd10;
        rom[520][7] = -8'd22;
        rom[520][8] = -8'd5;
        rom[520][9] = -8'd25;
        rom[520][10] = 8'd3;
        rom[520][11] = 8'd36;
        rom[520][12] = -8'd9;
        rom[520][13] = -8'd13;
        rom[520][14] = 8'd27;
        rom[520][15] = 8'd15;
        rom[520][16] = -8'd12;
        rom[520][17] = 8'd22;
        rom[520][18] = -8'd7;
        rom[520][19] = -8'd3;
        rom[520][20] = 8'd2;
        rom[520][21] = -8'd47;
        rom[520][22] = -8'd24;
        rom[520][23] = 8'd6;
        rom[520][24] = 8'd25;
        rom[520][25] = 8'd12;
        rom[520][26] = 8'd24;
        rom[520][27] = -8'd16;
        rom[520][28] = -8'd12;
        rom[520][29] = 8'd2;
        rom[520][30] = -8'd13;
        rom[520][31] = -8'd6;
        rom[520][32] = -8'd10;
        rom[520][33] = 8'd9;
        rom[520][34] = -8'd10;
        rom[520][35] = 8'd16;
        rom[520][36] = -8'd34;
        rom[520][37] = -8'd10;
        rom[520][38] = -8'd55;
        rom[520][39] = 8'd9;
        rom[520][40] = -8'd29;
        rom[520][41] = -8'd25;
        rom[520][42] = 8'd14;
        rom[520][43] = 8'd3;
        rom[520][44] = 8'd4;
        rom[520][45] = -8'd19;
        rom[520][46] = -8'd8;
        rom[520][47] = -8'd49;
        rom[520][48] = -8'd36;
        rom[520][49] = 8'd22;
        rom[520][50] = -8'd13;
        rom[520][51] = 8'd22;
        rom[520][52] = -8'd2;
        rom[520][53] = 8'd14;
        rom[520][54] = -8'd37;
        rom[520][55] = -8'd25;
        rom[520][56] = 8'd1;
        rom[520][57] = 8'd3;
        rom[520][58] = 8'd23;
        rom[520][59] = -8'd9;
        rom[520][60] = 8'd6;
        rom[520][61] = -8'd15;
        rom[520][62] = -8'd25;
        rom[520][63] = -8'd52;
        rom[521][0] = 8'd21;
        rom[521][1] = -8'd1;
        rom[521][2] = 8'd4;
        rom[521][3] = 8'd28;
        rom[521][4] = 8'd6;
        rom[521][5] = -8'd23;
        rom[521][6] = -8'd32;
        rom[521][7] = -8'd20;
        rom[521][8] = 8'd0;
        rom[521][9] = -8'd44;
        rom[521][10] = -8'd2;
        rom[521][11] = -8'd7;
        rom[521][12] = 8'd16;
        rom[521][13] = -8'd11;
        rom[521][14] = 8'd8;
        rom[521][15] = 8'd8;
        rom[521][16] = 8'd4;
        rom[521][17] = 8'd33;
        rom[521][18] = 8'd36;
        rom[521][19] = -8'd39;
        rom[521][20] = -8'd6;
        rom[521][21] = 8'd37;
        rom[521][22] = 8'd57;
        rom[521][23] = -8'd5;
        rom[521][24] = -8'd34;
        rom[521][25] = -8'd24;
        rom[521][26] = -8'd18;
        rom[521][27] = -8'd14;
        rom[521][28] = -8'd53;
        rom[521][29] = 8'd10;
        rom[521][30] = -8'd30;
        rom[521][31] = 8'd27;
        rom[521][32] = -8'd17;
        rom[521][33] = 8'd12;
        rom[521][34] = 8'd44;
        rom[521][35] = -8'd6;
        rom[521][36] = 8'd48;
        rom[521][37] = -8'd89;
        rom[521][38] = 8'd8;
        rom[521][39] = -8'd40;
        rom[521][40] = 8'd14;
        rom[521][41] = 8'd23;
        rom[521][42] = 8'd11;
        rom[521][43] = 8'd20;
        rom[521][44] = -8'd10;
        rom[521][45] = 8'd19;
        rom[521][46] = -8'd20;
        rom[521][47] = -8'd37;
        rom[521][48] = 8'd37;
        rom[521][49] = -8'd53;
        rom[521][50] = 8'd39;
        rom[521][51] = 8'd35;
        rom[521][52] = -8'd37;
        rom[521][53] = 8'd27;
        rom[521][54] = -8'd11;
        rom[521][55] = 8'd11;
        rom[521][56] = -8'd37;
        rom[521][57] = 8'd7;
        rom[521][58] = 8'd5;
        rom[521][59] = 8'd17;
        rom[521][60] = -8'd57;
        rom[521][61] = 8'd29;
        rom[521][62] = -8'd28;
        rom[521][63] = -8'd6;
        rom[522][0] = 8'd43;
        rom[522][1] = -8'd8;
        rom[522][2] = 8'd17;
        rom[522][3] = -8'd21;
        rom[522][4] = -8'd61;
        rom[522][5] = 8'd14;
        rom[522][6] = -8'd4;
        rom[522][7] = -8'd1;
        rom[522][8] = 8'd10;
        rom[522][9] = 8'd10;
        rom[522][10] = -8'd52;
        rom[522][11] = 8'd6;
        rom[522][12] = -8'd14;
        rom[522][13] = 8'd15;
        rom[522][14] = -8'd16;
        rom[522][15] = 8'd40;
        rom[522][16] = -8'd55;
        rom[522][17] = 8'd15;
        rom[522][18] = 8'd34;
        rom[522][19] = -8'd62;
        rom[522][20] = 8'd6;
        rom[522][21] = -8'd29;
        rom[522][22] = -8'd33;
        rom[522][23] = -8'd37;
        rom[522][24] = -8'd31;
        rom[522][25] = -8'd31;
        rom[522][26] = -8'd22;
        rom[522][27] = 8'd10;
        rom[522][28] = 8'd38;
        rom[522][29] = 8'd33;
        rom[522][30] = -8'd7;
        rom[522][31] = 8'd58;
        rom[522][32] = 8'd4;
        rom[522][33] = -8'd11;
        rom[522][34] = -8'd18;
        rom[522][35] = -8'd33;
        rom[522][36] = -8'd1;
        rom[522][37] = 8'd20;
        rom[522][38] = 8'd25;
        rom[522][39] = -8'd14;
        rom[522][40] = -8'd3;
        rom[522][41] = 8'd1;
        rom[522][42] = 8'd1;
        rom[522][43] = -8'd1;
        rom[522][44] = -8'd15;
        rom[522][45] = -8'd9;
        rom[522][46] = 8'd0;
        rom[522][47] = -8'd1;
        rom[522][48] = -8'd20;
        rom[522][49] = 8'd21;
        rom[522][50] = 8'd27;
        rom[522][51] = -8'd7;
        rom[522][52] = 8'd24;
        rom[522][53] = 8'd7;
        rom[522][54] = 8'd17;
        rom[522][55] = -8'd22;
        rom[522][56] = -8'd14;
        rom[522][57] = 8'd3;
        rom[522][58] = 8'd6;
        rom[522][59] = 8'd47;
        rom[522][60] = 8'd18;
        rom[522][61] = -8'd17;
        rom[522][62] = 8'd13;
        rom[522][63] = 8'd13;
        rom[523][0] = -8'd5;
        rom[523][1] = 8'd18;
        rom[523][2] = -8'd38;
        rom[523][3] = 8'd0;
        rom[523][4] = 8'd5;
        rom[523][5] = -8'd40;
        rom[523][6] = -8'd7;
        rom[523][7] = -8'd20;
        rom[523][8] = -8'd59;
        rom[523][9] = -8'd17;
        rom[523][10] = 8'd8;
        rom[523][11] = -8'd29;
        rom[523][12] = -8'd36;
        rom[523][13] = -8'd72;
        rom[523][14] = -8'd3;
        rom[523][15] = 8'd43;
        rom[523][16] = 8'd12;
        rom[523][17] = -8'd2;
        rom[523][18] = -8'd39;
        rom[523][19] = -8'd21;
        rom[523][20] = 8'd1;
        rom[523][21] = 8'd15;
        rom[523][22] = 8'd5;
        rom[523][23] = -8'd24;
        rom[523][24] = -8'd16;
        rom[523][25] = -8'd10;
        rom[523][26] = 8'd44;
        rom[523][27] = 8'd40;
        rom[523][28] = 8'd28;
        rom[523][29] = -8'd31;
        rom[523][30] = 8'd2;
        rom[523][31] = -8'd105;
        rom[523][32] = -8'd53;
        rom[523][33] = -8'd4;
        rom[523][34] = 8'd40;
        rom[523][35] = 8'd42;
        rom[523][36] = -8'd34;
        rom[523][37] = 8'd6;
        rom[523][38] = -8'd1;
        rom[523][39] = 8'd26;
        rom[523][40] = -8'd21;
        rom[523][41] = 8'd17;
        rom[523][42] = 8'd3;
        rom[523][43] = 8'd45;
        rom[523][44] = -8'd13;
        rom[523][45] = -8'd50;
        rom[523][46] = 8'd36;
        rom[523][47] = 8'd32;
        rom[523][48] = 8'd4;
        rom[523][49] = -8'd12;
        rom[523][50] = 8'd1;
        rom[523][51] = -8'd24;
        rom[523][52] = 8'd32;
        rom[523][53] = -8'd17;
        rom[523][54] = -8'd5;
        rom[523][55] = -8'd3;
        rom[523][56] = 8'd15;
        rom[523][57] = -8'd41;
        rom[523][58] = -8'd27;
        rom[523][59] = -8'd45;
        rom[523][60] = -8'd7;
        rom[523][61] = -8'd31;
        rom[523][62] = 8'd33;
        rom[523][63] = -8'd11;
        rom[524][0] = -8'd19;
        rom[524][1] = -8'd66;
        rom[524][2] = -8'd2;
        rom[524][3] = 8'd30;
        rom[524][4] = -8'd6;
        rom[524][5] = 8'd36;
        rom[524][6] = -8'd39;
        rom[524][7] = 8'd2;
        rom[524][8] = 8'd24;
        rom[524][9] = -8'd30;
        rom[524][10] = -8'd50;
        rom[524][11] = -8'd35;
        rom[524][12] = -8'd4;
        rom[524][13] = -8'd57;
        rom[524][14] = 8'd29;
        rom[524][15] = 8'd50;
        rom[524][16] = -8'd18;
        rom[524][17] = 8'd9;
        rom[524][18] = 8'd26;
        rom[524][19] = -8'd38;
        rom[524][20] = -8'd2;
        rom[524][21] = 8'd17;
        rom[524][22] = 8'd6;
        rom[524][23] = -8'd31;
        rom[524][24] = 8'd12;
        rom[524][25] = 8'd7;
        rom[524][26] = 8'd7;
        rom[524][27] = 8'd29;
        rom[524][28] = -8'd5;
        rom[524][29] = -8'd9;
        rom[524][30] = -8'd24;
        rom[524][31] = 8'd4;
        rom[524][32] = 8'd39;
        rom[524][33] = -8'd2;
        rom[524][34] = -8'd36;
        rom[524][35] = 8'd34;
        rom[524][36] = 8'd32;
        rom[524][37] = 8'd17;
        rom[524][38] = 8'd16;
        rom[524][39] = -8'd6;
        rom[524][40] = -8'd36;
        rom[524][41] = 8'd21;
        rom[524][42] = 8'd20;
        rom[524][43] = 8'd13;
        rom[524][44] = 8'd13;
        rom[524][45] = 8'd17;
        rom[524][46] = 8'd22;
        rom[524][47] = 8'd36;
        rom[524][48] = -8'd32;
        rom[524][49] = -8'd5;
        rom[524][50] = 8'd45;
        rom[524][51] = -8'd15;
        rom[524][52] = -8'd20;
        rom[524][53] = -8'd14;
        rom[524][54] = -8'd29;
        rom[524][55] = 8'd11;
        rom[524][56] = -8'd11;
        rom[524][57] = 8'd28;
        rom[524][58] = 8'd29;
        rom[524][59] = 8'd1;
        rom[524][60] = -8'd7;
        rom[524][61] = 8'd15;
        rom[524][62] = -8'd4;
        rom[524][63] = -8'd5;
        rom[525][0] = -8'd2;
        rom[525][1] = 8'd14;
        rom[525][2] = 8'd19;
        rom[525][3] = -8'd11;
        rom[525][4] = -8'd28;
        rom[525][5] = 8'd57;
        rom[525][6] = 8'd11;
        rom[525][7] = 8'd25;
        rom[525][8] = 8'd24;
        rom[525][9] = 8'd2;
        rom[525][10] = -8'd26;
        rom[525][11] = 8'd0;
        rom[525][12] = -8'd32;
        rom[525][13] = -8'd14;
        rom[525][14] = -8'd2;
        rom[525][15] = 8'd7;
        rom[525][16] = -8'd39;
        rom[525][17] = -8'd61;
        rom[525][18] = -8'd11;
        rom[525][19] = 8'd8;
        rom[525][20] = 8'd1;
        rom[525][21] = 8'd15;
        rom[525][22] = -8'd16;
        rom[525][23] = -8'd17;
        rom[525][24] = 8'd56;
        rom[525][25] = 8'd21;
        rom[525][26] = -8'd3;
        rom[525][27] = 8'd25;
        rom[525][28] = -8'd27;
        rom[525][29] = 8'd8;
        rom[525][30] = -8'd11;
        rom[525][31] = -8'd8;
        rom[525][32] = -8'd10;
        rom[525][33] = -8'd19;
        rom[525][34] = -8'd5;
        rom[525][35] = -8'd7;
        rom[525][36] = -8'd33;
        rom[525][37] = 8'd12;
        rom[525][38] = -8'd25;
        rom[525][39] = 8'd8;
        rom[525][40] = 8'd42;
        rom[525][41] = -8'd7;
        rom[525][42] = -8'd34;
        rom[525][43] = 8'd17;
        rom[525][44] = -8'd8;
        rom[525][45] = -8'd8;
        rom[525][46] = -8'd12;
        rom[525][47] = 8'd6;
        rom[525][48] = 8'd47;
        rom[525][49] = 8'd2;
        rom[525][50] = 8'd22;
        rom[525][51] = 8'd11;
        rom[525][52] = -8'd11;
        rom[525][53] = 8'd0;
        rom[525][54] = 8'd18;
        rom[525][55] = -8'd42;
        rom[525][56] = -8'd17;
        rom[525][57] = -8'd23;
        rom[525][58] = 8'd41;
        rom[525][59] = 8'd29;
        rom[525][60] = 8'd14;
        rom[525][61] = -8'd5;
        rom[525][62] = 8'd60;
        rom[525][63] = -8'd21;
        rom[526][0] = 8'd0;
        rom[526][1] = -8'd12;
        rom[526][2] = 8'd13;
        rom[526][3] = 8'd5;
        rom[526][4] = -8'd29;
        rom[526][5] = -8'd45;
        rom[526][6] = -8'd19;
        rom[526][7] = 8'd12;
        rom[526][8] = -8'd12;
        rom[526][9] = -8'd57;
        rom[526][10] = 8'd8;
        rom[526][11] = -8'd7;
        rom[526][12] = -8'd68;
        rom[526][13] = -8'd26;
        rom[526][14] = 8'd12;
        rom[526][15] = 8'd31;
        rom[526][16] = 8'd6;
        rom[526][17] = 8'd21;
        rom[526][18] = -8'd27;
        rom[526][19] = 8'd38;
        rom[526][20] = -8'd3;
        rom[526][21] = -8'd11;
        rom[526][22] = 8'd11;
        rom[526][23] = -8'd24;
        rom[526][24] = 8'd16;
        rom[526][25] = 8'd0;
        rom[526][26] = -8'd2;
        rom[526][27] = -8'd44;
        rom[526][28] = 8'd13;
        rom[526][29] = -8'd31;
        rom[526][30] = 8'd2;
        rom[526][31] = -8'd24;
        rom[526][32] = -8'd4;
        rom[526][33] = -8'd38;
        rom[526][34] = -8'd10;
        rom[526][35] = 8'd19;
        rom[526][36] = -8'd13;
        rom[526][37] = 8'd3;
        rom[526][38] = -8'd20;
        rom[526][39] = 8'd14;
        rom[526][40] = -8'd1;
        rom[526][41] = -8'd53;
        rom[526][42] = -8'd39;
        rom[526][43] = 8'd10;
        rom[526][44] = 8'd34;
        rom[526][45] = -8'd64;
        rom[526][46] = -8'd51;
        rom[526][47] = 8'd4;
        rom[526][48] = -8'd20;
        rom[526][49] = 8'd6;
        rom[526][50] = -8'd16;
        rom[526][51] = -8'd2;
        rom[526][52] = 8'd11;
        rom[526][53] = -8'd29;
        rom[526][54] = -8'd43;
        rom[526][55] = -8'd19;
        rom[526][56] = -8'd21;
        rom[526][57] = 8'd4;
        rom[526][58] = -8'd7;
        rom[526][59] = -8'd23;
        rom[526][60] = 8'd17;
        rom[526][61] = 8'd13;
        rom[526][62] = 8'd0;
        rom[526][63] = 8'd11;
        rom[527][0] = 8'd22;
        rom[527][1] = -8'd13;
        rom[527][2] = 8'd18;
        rom[527][3] = -8'd28;
        rom[527][4] = 8'd15;
        rom[527][5] = -8'd30;
        rom[527][6] = -8'd6;
        rom[527][7] = -8'd16;
        rom[527][8] = 8'd17;
        rom[527][9] = 8'd34;
        rom[527][10] = -8'd14;
        rom[527][11] = 8'd5;
        rom[527][12] = -8'd6;
        rom[527][13] = -8'd4;
        rom[527][14] = -8'd12;
        rom[527][15] = 8'd3;
        rom[527][16] = 8'd0;
        rom[527][17] = 8'd22;
        rom[527][18] = 8'd23;
        rom[527][19] = -8'd37;
        rom[527][20] = -8'd4;
        rom[527][21] = -8'd19;
        rom[527][22] = 8'd1;
        rom[527][23] = -8'd31;
        rom[527][24] = 8'd7;
        rom[527][25] = -8'd14;
        rom[527][26] = 8'd3;
        rom[527][27] = -8'd47;
        rom[527][28] = -8'd3;
        rom[527][29] = -8'd8;
        rom[527][30] = 8'd11;
        rom[527][31] = 8'd48;
        rom[527][32] = -8'd20;
        rom[527][33] = -8'd10;
        rom[527][34] = -8'd34;
        rom[527][35] = -8'd14;
        rom[527][36] = -8'd14;
        rom[527][37] = -8'd75;
        rom[527][38] = 8'd0;
        rom[527][39] = 8'd12;
        rom[527][40] = 8'd63;
        rom[527][41] = -8'd28;
        rom[527][42] = 8'd1;
        rom[527][43] = 8'd8;
        rom[527][44] = 8'd37;
        rom[527][45] = -8'd33;
        rom[527][46] = -8'd34;
        rom[527][47] = -8'd25;
        rom[527][48] = 8'd21;
        rom[527][49] = -8'd3;
        rom[527][50] = -8'd4;
        rom[527][51] = 8'd36;
        rom[527][52] = 8'd5;
        rom[527][53] = 8'd8;
        rom[527][54] = -8'd17;
        rom[527][55] = -8'd8;
        rom[527][56] = -8'd9;
        rom[527][57] = 8'd21;
        rom[527][58] = -8'd32;
        rom[527][59] = -8'd26;
        rom[527][60] = 8'd20;
        rom[527][61] = -8'd44;
        rom[527][62] = -8'd6;
        rom[527][63] = -8'd23;
        rom[528][0] = -8'd1;
        rom[528][1] = 8'd1;
        rom[528][2] = 8'd9;
        rom[528][3] = -8'd5;
        rom[528][4] = -8'd3;
        rom[528][5] = -8'd3;
        rom[528][6] = 8'd6;
        rom[528][7] = -8'd5;
        rom[528][8] = -8'd8;
        rom[528][9] = 8'd1;
        rom[528][10] = -8'd3;
        rom[528][11] = -8'd6;
        rom[528][12] = 8'd1;
        rom[528][13] = 8'd3;
        rom[528][14] = -8'd5;
        rom[528][15] = 8'd0;
        rom[528][16] = 8'd6;
        rom[528][17] = -8'd5;
        rom[528][18] = 8'd2;
        rom[528][19] = -8'd6;
        rom[528][20] = -8'd2;
        rom[528][21] = -8'd2;
        rom[528][22] = -8'd1;
        rom[528][23] = 8'd2;
        rom[528][24] = -8'd2;
        rom[528][25] = -8'd4;
        rom[528][26] = 8'd3;
        rom[528][27] = -8'd1;
        rom[528][28] = -8'd2;
        rom[528][29] = -8'd8;
        rom[528][30] = 8'd4;
        rom[528][31] = -8'd2;
        rom[528][32] = 8'd3;
        rom[528][33] = -8'd7;
        rom[528][34] = 8'd1;
        rom[528][35] = -8'd4;
        rom[528][36] = 8'd8;
        rom[528][37] = 8'd6;
        rom[528][38] = 8'd7;
        rom[528][39] = -8'd9;
        rom[528][40] = -8'd2;
        rom[528][41] = 8'd2;
        rom[528][42] = 8'd8;
        rom[528][43] = 8'd0;
        rom[528][44] = 8'd9;
        rom[528][45] = -8'd4;
        rom[528][46] = -8'd5;
        rom[528][47] = 8'd1;
        rom[528][48] = 8'd6;
        rom[528][49] = -8'd4;
        rom[528][50] = -8'd7;
        rom[528][51] = 8'd1;
        rom[528][52] = 8'd9;
        rom[528][53] = -8'd8;
        rom[528][54] = 8'd3;
        rom[528][55] = -8'd1;
        rom[528][56] = 8'd3;
        rom[528][57] = 8'd5;
        rom[528][58] = 8'd5;
        rom[528][59] = -8'd7;
        rom[528][60] = 8'd5;
        rom[528][61] = -8'd9;
        rom[528][62] = -8'd7;
        rom[528][63] = -8'd7;
        rom[529][0] = 8'd25;
        rom[529][1] = -8'd6;
        rom[529][2] = -8'd58;
        rom[529][3] = 8'd8;
        rom[529][4] = 8'd27;
        rom[529][5] = -8'd21;
        rom[529][6] = 8'd26;
        rom[529][7] = -8'd17;
        rom[529][8] = -8'd40;
        rom[529][9] = 8'd4;
        rom[529][10] = -8'd53;
        rom[529][11] = 8'd11;
        rom[529][12] = -8'd22;
        rom[529][13] = 8'd14;
        rom[529][14] = 8'd5;
        rom[529][15] = -8'd15;
        rom[529][16] = 8'd24;
        rom[529][17] = 8'd9;
        rom[529][18] = 8'd2;
        rom[529][19] = -8'd71;
        rom[529][20] = -8'd12;
        rom[529][21] = 8'd22;
        rom[529][22] = 8'd12;
        rom[529][23] = -8'd7;
        rom[529][24] = 8'd26;
        rom[529][25] = 8'd14;
        rom[529][26] = -8'd18;
        rom[529][27] = 8'd37;
        rom[529][28] = -8'd15;
        rom[529][29] = -8'd27;
        rom[529][30] = -8'd9;
        rom[529][31] = -8'd8;
        rom[529][32] = -8'd21;
        rom[529][33] = 8'd7;
        rom[529][34] = -8'd45;
        rom[529][35] = 8'd14;
        rom[529][36] = 8'd36;
        rom[529][37] = 8'd15;
        rom[529][38] = 8'd1;
        rom[529][39] = 8'd17;
        rom[529][40] = -8'd10;
        rom[529][41] = -8'd17;
        rom[529][42] = -8'd53;
        rom[529][43] = 8'd23;
        rom[529][44] = -8'd8;
        rom[529][45] = 8'd36;
        rom[529][46] = 8'd3;
        rom[529][47] = -8'd20;
        rom[529][48] = 8'd27;
        rom[529][49] = 8'd17;
        rom[529][50] = 8'd3;
        rom[529][51] = 8'd9;
        rom[529][52] = 8'd39;
        rom[529][53] = 8'd20;
        rom[529][54] = -8'd30;
        rom[529][55] = 8'd27;
        rom[529][56] = -8'd11;
        rom[529][57] = -8'd29;
        rom[529][58] = -8'd45;
        rom[529][59] = 8'd10;
        rom[529][60] = 8'd31;
        rom[529][61] = 8'd37;
        rom[529][62] = 8'd18;
        rom[529][63] = -8'd22;
        rom[530][0] = 8'd11;
        rom[530][1] = -8'd16;
        rom[530][2] = 8'd4;
        rom[530][3] = -8'd51;
        rom[530][4] = -8'd14;
        rom[530][5] = 8'd20;
        rom[530][6] = 8'd18;
        rom[530][7] = -8'd24;
        rom[530][8] = 8'd16;
        rom[530][9] = -8'd25;
        rom[530][10] = -8'd61;
        rom[530][11] = 8'd11;
        rom[530][12] = -8'd23;
        rom[530][13] = -8'd25;
        rom[530][14] = 8'd2;
        rom[530][15] = 8'd12;
        rom[530][16] = -8'd81;
        rom[530][17] = -8'd47;
        rom[530][18] = -8'd25;
        rom[530][19] = -8'd16;
        rom[530][20] = 8'd2;
        rom[530][21] = -8'd11;
        rom[530][22] = 8'd3;
        rom[530][23] = -8'd5;
        rom[530][24] = -8'd16;
        rom[530][25] = -8'd12;
        rom[530][26] = 8'd16;
        rom[530][27] = 8'd6;
        rom[530][28] = -8'd44;
        rom[530][29] = -8'd26;
        rom[530][30] = 8'd29;
        rom[530][31] = -8'd14;
        rom[530][32] = 8'd2;
        rom[530][33] = -8'd25;
        rom[530][34] = -8'd1;
        rom[530][35] = -8'd19;
        rom[530][36] = -8'd8;
        rom[530][37] = -8'd22;
        rom[530][38] = -8'd23;
        rom[530][39] = 8'd4;
        rom[530][40] = -8'd27;
        rom[530][41] = 8'd26;
        rom[530][42] = -8'd9;
        rom[530][43] = 8'd40;
        rom[530][44] = 8'd7;
        rom[530][45] = -8'd79;
        rom[530][46] = -8'd21;
        rom[530][47] = -8'd65;
        rom[530][48] = 8'd22;
        rom[530][49] = -8'd8;
        rom[530][50] = -8'd4;
        rom[530][51] = -8'd1;
        rom[530][52] = 8'd5;
        rom[530][53] = 8'd28;
        rom[530][54] = 8'd4;
        rom[530][55] = 8'd12;
        rom[530][56] = -8'd18;
        rom[530][57] = 8'd4;
        rom[530][58] = -8'd36;
        rom[530][59] = -8'd33;
        rom[530][60] = -8'd25;
        rom[530][61] = -8'd24;
        rom[530][62] = -8'd26;
        rom[530][63] = -8'd9;
        rom[531][0] = 8'd26;
        rom[531][1] = 8'd8;
        rom[531][2] = 8'd15;
        rom[531][3] = -8'd24;
        rom[531][4] = 8'd8;
        rom[531][5] = -8'd22;
        rom[531][6] = -8'd3;
        rom[531][7] = 8'd8;
        rom[531][8] = -8'd28;
        rom[531][9] = -8'd3;
        rom[531][10] = -8'd50;
        rom[531][11] = -8'd20;
        rom[531][12] = 8'd10;
        rom[531][13] = 8'd35;
        rom[531][14] = 8'd32;
        rom[531][15] = 8'd35;
        rom[531][16] = 8'd39;
        rom[531][17] = 8'd12;
        rom[531][18] = -8'd12;
        rom[531][19] = 8'd23;
        rom[531][20] = 8'd3;
        rom[531][21] = -8'd20;
        rom[531][22] = 8'd5;
        rom[531][23] = 8'd13;
        rom[531][24] = 8'd19;
        rom[531][25] = -8'd31;
        rom[531][26] = 8'd3;
        rom[531][27] = -8'd7;
        rom[531][28] = -8'd9;
        rom[531][29] = 8'd18;
        rom[531][30] = -8'd10;
        rom[531][31] = -8'd44;
        rom[531][32] = 8'd37;
        rom[531][33] = 8'd3;
        rom[531][34] = 8'd18;
        rom[531][35] = -8'd77;
        rom[531][36] = 8'd33;
        rom[531][37] = -8'd69;
        rom[531][38] = -8'd4;
        rom[531][39] = -8'd7;
        rom[531][40] = -8'd12;
        rom[531][41] = -8'd22;
        rom[531][42] = 8'd7;
        rom[531][43] = -8'd12;
        rom[531][44] = 8'd21;
        rom[531][45] = 8'd1;
        rom[531][46] = 8'd14;
        rom[531][47] = -8'd10;
        rom[531][48] = 8'd21;
        rom[531][49] = -8'd33;
        rom[531][50] = -8'd12;
        rom[531][51] = 8'd7;
        rom[531][52] = 8'd24;
        rom[531][53] = 8'd14;
        rom[531][54] = -8'd12;
        rom[531][55] = 8'd1;
        rom[531][56] = -8'd32;
        rom[531][57] = 8'd41;
        rom[531][58] = -8'd35;
        rom[531][59] = 8'd3;
        rom[531][60] = 8'd9;
        rom[531][61] = 8'd3;
        rom[531][62] = 8'd5;
        rom[531][63] = -8'd13;
        rom[532][0] = 8'd10;
        rom[532][1] = 8'd35;
        rom[532][2] = -8'd40;
        rom[532][3] = 8'd4;
        rom[532][4] = -8'd100;
        rom[532][5] = 8'd23;
        rom[532][6] = -8'd17;
        rom[532][7] = -8'd10;
        rom[532][8] = -8'd22;
        rom[532][9] = -8'd15;
        rom[532][10] = -8'd8;
        rom[532][11] = 8'd38;
        rom[532][12] = 8'd8;
        rom[532][13] = 8'd15;
        rom[532][14] = -8'd34;
        rom[532][15] = 8'd6;
        rom[532][16] = -8'd19;
        rom[532][17] = 8'd3;
        rom[532][18] = 8'd14;
        rom[532][19] = 8'd14;
        rom[532][20] = -8'd14;
        rom[532][21] = 8'd0;
        rom[532][22] = 8'd10;
        rom[532][23] = 8'd25;
        rom[532][24] = 8'd15;
        rom[532][25] = 8'd0;
        rom[532][26] = -8'd12;
        rom[532][27] = -8'd18;
        rom[532][28] = -8'd27;
        rom[532][29] = -8'd40;
        rom[532][30] = -8'd22;
        rom[532][31] = -8'd44;
        rom[532][32] = -8'd30;
        rom[532][33] = -8'd26;
        rom[532][34] = 8'd8;
        rom[532][35] = -8'd32;
        rom[532][36] = -8'd5;
        rom[532][37] = -8'd4;
        rom[532][38] = 8'd38;
        rom[532][39] = -8'd15;
        rom[532][40] = 8'd38;
        rom[532][41] = -8'd10;
        rom[532][42] = 8'd42;
        rom[532][43] = -8'd26;
        rom[532][44] = 8'd2;
        rom[532][45] = -8'd28;
        rom[532][46] = 8'd3;
        rom[532][47] = 8'd21;
        rom[532][48] = 8'd0;
        rom[532][49] = 8'd22;
        rom[532][50] = -8'd58;
        rom[532][51] = -8'd16;
        rom[532][52] = 8'd8;
        rom[532][53] = -8'd43;
        rom[532][54] = -8'd4;
        rom[532][55] = 8'd9;
        rom[532][56] = -8'd14;
        rom[532][57] = 8'd0;
        rom[532][58] = 8'd12;
        rom[532][59] = -8'd20;
        rom[532][60] = 8'd21;
        rom[532][61] = -8'd12;
        rom[532][62] = -8'd36;
        rom[532][63] = -8'd3;
        rom[533][0] = 8'd3;
        rom[533][1] = -8'd9;
        rom[533][2] = 8'd2;
        rom[533][3] = 8'd1;
        rom[533][4] = 8'd4;
        rom[533][5] = -8'd2;
        rom[533][6] = -8'd7;
        rom[533][7] = 8'd5;
        rom[533][8] = 8'd6;
        rom[533][9] = -8'd6;
        rom[533][10] = -8'd3;
        rom[533][11] = 8'd1;
        rom[533][12] = 8'd0;
        rom[533][13] = -8'd1;
        rom[533][14] = 8'd5;
        rom[533][15] = -8'd6;
        rom[533][16] = 8'd8;
        rom[533][17] = -8'd1;
        rom[533][18] = 8'd1;
        rom[533][19] = 8'd0;
        rom[533][20] = -8'd7;
        rom[533][21] = 8'd0;
        rom[533][22] = 8'd6;
        rom[533][23] = -8'd3;
        rom[533][24] = 8'd1;
        rom[533][25] = 8'd0;
        rom[533][26] = -8'd6;
        rom[533][27] = -8'd8;
        rom[533][28] = 8'd6;
        rom[533][29] = 8'd9;
        rom[533][30] = -8'd6;
        rom[533][31] = 8'd1;
        rom[533][32] = -8'd6;
        rom[533][33] = -8'd5;
        rom[533][34] = -8'd1;
        rom[533][35] = 8'd0;
        rom[533][36] = 8'd9;
        rom[533][37] = 8'd0;
        rom[533][38] = 8'd8;
        rom[533][39] = -8'd6;
        rom[533][40] = 8'd6;
        rom[533][41] = -8'd6;
        rom[533][42] = 8'd3;
        rom[533][43] = -8'd4;
        rom[533][44] = 8'd12;
        rom[533][45] = 8'd0;
        rom[533][46] = 8'd4;
        rom[533][47] = -8'd9;
        rom[533][48] = 8'd9;
        rom[533][49] = -8'd1;
        rom[533][50] = 8'd2;
        rom[533][51] = -8'd2;
        rom[533][52] = 8'd2;
        rom[533][53] = -8'd3;
        rom[533][54] = -8'd9;
        rom[533][55] = 8'd7;
        rom[533][56] = -8'd1;
        rom[533][57] = -8'd3;
        rom[533][58] = -8'd5;
        rom[533][59] = -8'd9;
        rom[533][60] = 8'd7;
        rom[533][61] = -8'd5;
        rom[533][62] = -8'd4;
        rom[533][63] = -8'd5;
        rom[534][0] = -8'd47;
        rom[534][1] = 8'd45;
        rom[534][2] = -8'd16;
        rom[534][3] = 8'd1;
        rom[534][4] = 8'd2;
        rom[534][5] = -8'd56;
        rom[534][6] = -8'd10;
        rom[534][7] = -8'd93;
        rom[534][8] = 8'd1;
        rom[534][9] = 8'd32;
        rom[534][10] = -8'd49;
        rom[534][11] = -8'd3;
        rom[534][12] = -8'd16;
        rom[534][13] = -8'd101;
        rom[534][14] = -8'd8;
        rom[534][15] = -8'd9;
        rom[534][16] = 8'd6;
        rom[534][17] = 8'd17;
        rom[534][18] = -8'd23;
        rom[534][19] = 8'd42;
        rom[534][20] = 8'd4;
        rom[534][21] = 8'd13;
        rom[534][22] = -8'd57;
        rom[534][23] = 8'd10;
        rom[534][24] = -8'd15;
        rom[534][25] = 8'd33;
        rom[534][26] = -8'd5;
        rom[534][27] = 8'd20;
        rom[534][28] = -8'd7;
        rom[534][29] = 8'd39;
        rom[534][30] = -8'd15;
        rom[534][31] = 8'd10;
        rom[534][32] = -8'd37;
        rom[534][33] = 8'd11;
        rom[534][34] = 8'd31;
        rom[534][35] = -8'd40;
        rom[534][36] = 8'd0;
        rom[534][37] = 8'd23;
        rom[534][38] = 8'd30;
        rom[534][39] = 8'd11;
        rom[534][40] = -8'd31;
        rom[534][41] = 8'd34;
        rom[534][42] = 8'd16;
        rom[534][43] = 8'd30;
        rom[534][44] = -8'd35;
        rom[534][45] = 8'd30;
        rom[534][46] = -8'd36;
        rom[534][47] = 8'd19;
        rom[534][48] = -8'd8;
        rom[534][49] = -8'd2;
        rom[534][50] = 8'd23;
        rom[534][51] = -8'd3;
        rom[534][52] = 8'd28;
        rom[534][53] = 8'd14;
        rom[534][54] = 8'd38;
        rom[534][55] = -8'd7;
        rom[534][56] = -8'd40;
        rom[534][57] = 8'd7;
        rom[534][58] = 8'd23;
        rom[534][59] = 8'd27;
        rom[534][60] = -8'd5;
        rom[534][61] = -8'd9;
        rom[534][62] = -8'd11;
        rom[534][63] = 8'd33;
        rom[535][0] = -8'd16;
        rom[535][1] = 8'd20;
        rom[535][2] = -8'd12;
        rom[535][3] = 8'd13;
        rom[535][4] = 8'd10;
        rom[535][5] = 8'd14;
        rom[535][6] = -8'd25;
        rom[535][7] = -8'd10;
        rom[535][8] = -8'd50;
        rom[535][9] = 8'd19;
        rom[535][10] = -8'd21;
        rom[535][11] = 8'd28;
        rom[535][12] = 8'd4;
        rom[535][13] = -8'd6;
        rom[535][14] = -8'd34;
        rom[535][15] = -8'd45;
        rom[535][16] = -8'd52;
        rom[535][17] = -8'd48;
        rom[535][18] = -8'd21;
        rom[535][19] = -8'd15;
        rom[535][20] = -8'd12;
        rom[535][21] = 8'd7;
        rom[535][22] = -8'd19;
        rom[535][23] = -8'd23;
        rom[535][24] = 8'd45;
        rom[535][25] = -8'd28;
        rom[535][26] = -8'd37;
        rom[535][27] = 8'd7;
        rom[535][28] = 8'd5;
        rom[535][29] = -8'd4;
        rom[535][30] = 8'd15;
        rom[535][31] = -8'd36;
        rom[535][32] = -8'd2;
        rom[535][33] = -8'd28;
        rom[535][34] = 8'd32;
        rom[535][35] = 8'd26;
        rom[535][36] = -8'd8;
        rom[535][37] = -8'd7;
        rom[535][38] = -8'd3;
        rom[535][39] = -8'd2;
        rom[535][40] = -8'd4;
        rom[535][41] = -8'd23;
        rom[535][42] = -8'd11;
        rom[535][43] = -8'd4;
        rom[535][44] = 8'd10;
        rom[535][45] = -8'd45;
        rom[535][46] = -8'd12;
        rom[535][47] = 8'd62;
        rom[535][48] = -8'd35;
        rom[535][49] = 8'd34;
        rom[535][50] = -8'd26;
        rom[535][51] = -8'd17;
        rom[535][52] = -8'd16;
        rom[535][53] = -8'd7;
        rom[535][54] = -8'd43;
        rom[535][55] = -8'd5;
        rom[535][56] = 8'd2;
        rom[535][57] = -8'd12;
        rom[535][58] = 8'd16;
        rom[535][59] = 8'd17;
        rom[535][60] = 8'd7;
        rom[535][61] = 8'd2;
        rom[535][62] = -8'd15;
        rom[535][63] = -8'd13;
        rom[536][0] = -8'd32;
        rom[536][1] = -8'd39;
        rom[536][2] = -8'd2;
        rom[536][3] = 8'd29;
        rom[536][4] = 8'd21;
        rom[536][5] = -8'd12;
        rom[536][6] = -8'd6;
        rom[536][7] = 8'd34;
        rom[536][8] = -8'd40;
        rom[536][9] = -8'd10;
        rom[536][10] = -8'd18;
        rom[536][11] = 8'd7;
        rom[536][12] = 8'd15;
        rom[536][13] = 8'd13;
        rom[536][14] = -8'd21;
        rom[536][15] = 8'd17;
        rom[536][16] = 8'd32;
        rom[536][17] = 8'd5;
        rom[536][18] = 8'd1;
        rom[536][19] = 8'd33;
        rom[536][20] = -8'd7;
        rom[536][21] = -8'd5;
        rom[536][22] = 8'd10;
        rom[536][23] = -8'd39;
        rom[536][24] = 8'd18;
        rom[536][25] = -8'd53;
        rom[536][26] = 8'd45;
        rom[536][27] = 8'd32;
        rom[536][28] = -8'd4;
        rom[536][29] = 8'd1;
        rom[536][30] = 8'd4;
        rom[536][31] = -8'd1;
        rom[536][32] = 8'd37;
        rom[536][33] = 8'd54;
        rom[536][34] = -8'd18;
        rom[536][35] = 8'd25;
        rom[536][36] = 8'd25;
        rom[536][37] = 8'd22;
        rom[536][38] = -8'd21;
        rom[536][39] = 8'd16;
        rom[536][40] = 8'd36;
        rom[536][41] = -8'd4;
        rom[536][42] = 8'd9;
        rom[536][43] = 8'd2;
        rom[536][44] = -8'd32;
        rom[536][45] = 8'd19;
        rom[536][46] = 8'd21;
        rom[536][47] = -8'd2;
        rom[536][48] = -8'd46;
        rom[536][49] = 8'd4;
        rom[536][50] = 8'd12;
        rom[536][51] = -8'd29;
        rom[536][52] = 8'd20;
        rom[536][53] = -8'd1;
        rom[536][54] = 8'd7;
        rom[536][55] = -8'd45;
        rom[536][56] = 8'd4;
        rom[536][57] = -8'd9;
        rom[536][58] = -8'd3;
        rom[536][59] = 8'd11;
        rom[536][60] = 8'd14;
        rom[536][61] = 8'd13;
        rom[536][62] = 8'd37;
        rom[536][63] = 8'd11;
        rom[537][0] = 8'd28;
        rom[537][1] = 8'd0;
        rom[537][2] = -8'd53;
        rom[537][3] = -8'd24;
        rom[537][4] = -8'd4;
        rom[537][5] = -8'd9;
        rom[537][6] = 8'd32;
        rom[537][7] = 8'd16;
        rom[537][8] = -8'd16;
        rom[537][9] = 8'd0;
        rom[537][10] = -8'd20;
        rom[537][11] = -8'd16;
        rom[537][12] = 8'd9;
        rom[537][13] = -8'd70;
        rom[537][14] = -8'd7;
        rom[537][15] = 8'd22;
        rom[537][16] = -8'd21;
        rom[537][17] = 8'd37;
        rom[537][18] = -8'd3;
        rom[537][19] = 8'd31;
        rom[537][20] = 8'd1;
        rom[537][21] = 8'd23;
        rom[537][22] = 8'd11;
        rom[537][23] = 8'd14;
        rom[537][24] = -8'd9;
        rom[537][25] = -8'd54;
        rom[537][26] = 8'd9;
        rom[537][27] = 8'd10;
        rom[537][28] = 8'd5;
        rom[537][29] = -8'd9;
        rom[537][30] = 8'd2;
        rom[537][31] = -8'd47;
        rom[537][32] = 8'd30;
        rom[537][33] = -8'd12;
        rom[537][34] = 8'd29;
        rom[537][35] = -8'd28;
        rom[537][36] = -8'd39;
        rom[537][37] = -8'd79;
        rom[537][38] = -8'd24;
        rom[537][39] = 8'd4;
        rom[537][40] = -8'd37;
        rom[537][41] = 8'd18;
        rom[537][42] = -8'd74;
        rom[537][43] = -8'd34;
        rom[537][44] = -8'd45;
        rom[537][45] = -8'd5;
        rom[537][46] = -8'd20;
        rom[537][47] = -8'd26;
        rom[537][48] = 8'd26;
        rom[537][49] = -8'd25;
        rom[537][50] = -8'd36;
        rom[537][51] = -8'd28;
        rom[537][52] = -8'd50;
        rom[537][53] = -8'd15;
        rom[537][54] = 8'd12;
        rom[537][55] = -8'd10;
        rom[537][56] = -8'd17;
        rom[537][57] = -8'd57;
        rom[537][58] = 8'd32;
        rom[537][59] = 8'd24;
        rom[537][60] = 8'd9;
        rom[537][61] = -8'd18;
        rom[537][62] = -8'd47;
        rom[537][63] = 8'd28;
        rom[538][0] = -8'd16;
        rom[538][1] = 8'd21;
        rom[538][2] = -8'd24;
        rom[538][3] = 8'd10;
        rom[538][4] = 8'd15;
        rom[538][5] = 8'd8;
        rom[538][6] = 8'd44;
        rom[538][7] = -8'd109;
        rom[538][8] = 8'd0;
        rom[538][9] = -8'd5;
        rom[538][10] = 8'd2;
        rom[538][11] = -8'd23;
        rom[538][12] = 8'd44;
        rom[538][13] = -8'd2;
        rom[538][14] = -8'd27;
        rom[538][15] = -8'd59;
        rom[538][16] = -8'd11;
        rom[538][17] = -8'd11;
        rom[538][18] = -8'd43;
        rom[538][19] = 8'd0;
        rom[538][20] = -8'd11;
        rom[538][21] = 8'd44;
        rom[538][22] = 8'd26;
        rom[538][23] = -8'd16;
        rom[538][24] = 8'd13;
        rom[538][25] = -8'd14;
        rom[538][26] = -8'd38;
        rom[538][27] = 8'd25;
        rom[538][28] = 8'd1;
        rom[538][29] = 8'd20;
        rom[538][30] = -8'd12;
        rom[538][31] = -8'd24;
        rom[538][32] = 8'd10;
        rom[538][33] = -8'd44;
        rom[538][34] = 8'd8;
        rom[538][35] = 8'd23;
        rom[538][36] = 8'd3;
        rom[538][37] = -8'd16;
        rom[538][38] = -8'd28;
        rom[538][39] = -8'd3;
        rom[538][40] = -8'd51;
        rom[538][41] = 8'd17;
        rom[538][42] = -8'd2;
        rom[538][43] = -8'd8;
        rom[538][44] = 8'd7;
        rom[538][45] = -8'd5;
        rom[538][46] = -8'd43;
        rom[538][47] = 8'd31;
        rom[538][48] = 8'd6;
        rom[538][49] = 8'd39;
        rom[538][50] = -8'd37;
        rom[538][51] = 8'd18;
        rom[538][52] = -8'd28;
        rom[538][53] = 8'd3;
        rom[538][54] = 8'd22;
        rom[538][55] = -8'd5;
        rom[538][56] = 8'd2;
        rom[538][57] = 8'd10;
        rom[538][58] = 8'd2;
        rom[538][59] = 8'd2;
        rom[538][60] = 8'd55;
        rom[538][61] = -8'd36;
        rom[538][62] = 8'd2;
        rom[538][63] = 8'd19;
        rom[539][0] = 8'd3;
        rom[539][1] = 8'd67;
        rom[539][2] = -8'd25;
        rom[539][3] = 8'd10;
        rom[539][4] = 8'd8;
        rom[539][5] = 8'd35;
        rom[539][6] = 8'd1;
        rom[539][7] = -8'd6;
        rom[539][8] = 8'd21;
        rom[539][9] = 8'd24;
        rom[539][10] = 8'd14;
        rom[539][11] = 8'd35;
        rom[539][12] = -8'd5;
        rom[539][13] = -8'd28;
        rom[539][14] = 8'd11;
        rom[539][15] = 8'd13;
        rom[539][16] = -8'd1;
        rom[539][17] = -8'd8;
        rom[539][18] = 8'd2;
        rom[539][19] = 8'd31;
        rom[539][20] = -8'd1;
        rom[539][21] = 8'd34;
        rom[539][22] = -8'd17;
        rom[539][23] = 8'd1;
        rom[539][24] = 8'd10;
        rom[539][25] = -8'd1;
        rom[539][26] = -8'd19;
        rom[539][27] = -8'd29;
        rom[539][28] = -8'd18;
        rom[539][29] = 8'd29;
        rom[539][30] = -8'd20;
        rom[539][31] = 8'd27;
        rom[539][32] = -8'd16;
        rom[539][33] = -8'd11;
        rom[539][34] = 8'd3;
        rom[539][35] = -8'd41;
        rom[539][36] = -8'd14;
        rom[539][37] = -8'd67;
        rom[539][38] = -8'd18;
        rom[539][39] = -8'd31;
        rom[539][40] = 8'd2;
        rom[539][41] = -8'd3;
        rom[539][42] = 8'd42;
        rom[539][43] = -8'd33;
        rom[539][44] = 8'd33;
        rom[539][45] = -8'd3;
        rom[539][46] = 8'd62;
        rom[539][47] = -8'd29;
        rom[539][48] = 8'd49;
        rom[539][49] = -8'd23;
        rom[539][50] = -8'd16;
        rom[539][51] = 8'd2;
        rom[539][52] = 8'd23;
        rom[539][53] = -8'd25;
        rom[539][54] = 8'd19;
        rom[539][55] = 8'd6;
        rom[539][56] = 8'd36;
        rom[539][57] = -8'd47;
        rom[539][58] = 8'd18;
        rom[539][59] = 8'd12;
        rom[539][60] = -8'd5;
        rom[539][61] = 8'd11;
        rom[539][62] = 8'd12;
        rom[539][63] = -8'd24;
        rom[540][0] = 8'd18;
        rom[540][1] = -8'd4;
        rom[540][2] = -8'd1;
        rom[540][3] = -8'd5;
        rom[540][4] = 8'd19;
        rom[540][5] = -8'd5;
        rom[540][6] = 8'd1;
        rom[540][7] = 8'd16;
        rom[540][8] = -8'd23;
        rom[540][9] = 8'd27;
        rom[540][10] = 8'd3;
        rom[540][11] = 8'd8;
        rom[540][12] = 8'd5;
        rom[540][13] = 8'd11;
        rom[540][14] = 8'd22;
        rom[540][15] = 8'd30;
        rom[540][16] = 8'd12;
        rom[540][17] = 8'd11;
        rom[540][18] = -8'd48;
        rom[540][19] = -8'd19;
        rom[540][20] = -8'd7;
        rom[540][21] = 8'd6;
        rom[540][22] = 8'd32;
        rom[540][23] = -8'd13;
        rom[540][24] = 8'd8;
        rom[540][25] = -8'd5;
        rom[540][26] = -8'd5;
        rom[540][27] = -8'd76;
        rom[540][28] = 8'd22;
        rom[540][29] = 8'd21;
        rom[540][30] = 8'd20;
        rom[540][31] = 8'd25;
        rom[540][32] = -8'd9;
        rom[540][33] = -8'd7;
        rom[540][34] = -8'd7;
        rom[540][35] = -8'd8;
        rom[540][36] = 8'd22;
        rom[540][37] = -8'd9;
        rom[540][38] = 8'd41;
        rom[540][39] = -8'd43;
        rom[540][40] = -8'd50;
        rom[540][41] = 8'd33;
        rom[540][42] = -8'd30;
        rom[540][43] = 8'd32;
        rom[540][44] = 8'd9;
        rom[540][45] = 8'd39;
        rom[540][46] = -8'd6;
        rom[540][47] = -8'd5;
        rom[540][48] = -8'd10;
        rom[540][49] = -8'd9;
        rom[540][50] = 8'd8;
        rom[540][51] = -8'd21;
        rom[540][52] = 8'd24;
        rom[540][53] = -8'd18;
        rom[540][54] = 8'd6;
        rom[540][55] = 8'd28;
        rom[540][56] = 8'd9;
        rom[540][57] = 8'd17;
        rom[540][58] = -8'd9;
        rom[540][59] = 8'd44;
        rom[540][60] = -8'd16;
        rom[540][61] = -8'd3;
        rom[540][62] = 8'd45;
        rom[540][63] = -8'd19;
        rom[541][0] = 8'd20;
        rom[541][1] = 8'd10;
        rom[541][2] = -8'd4;
        rom[541][3] = -8'd4;
        rom[541][4] = -8'd22;
        rom[541][5] = -8'd12;
        rom[541][6] = -8'd7;
        rom[541][7] = 8'd31;
        rom[541][8] = 8'd9;
        rom[541][9] = 8'd8;
        rom[541][10] = -8'd40;
        rom[541][11] = -8'd44;
        rom[541][12] = -8'd15;
        rom[541][13] = 8'd28;
        rom[541][14] = -8'd15;
        rom[541][15] = 8'd47;
        rom[541][16] = 8'd32;
        rom[541][17] = -8'd17;
        rom[541][18] = -8'd29;
        rom[541][19] = 8'd7;
        rom[541][20] = -8'd3;
        rom[541][21] = 8'd15;
        rom[541][22] = -8'd35;
        rom[541][23] = -8'd6;
        rom[541][24] = 8'd7;
        rom[541][25] = 8'd25;
        rom[541][26] = 8'd10;
        rom[541][27] = -8'd51;
        rom[541][28] = 8'd15;
        rom[541][29] = 8'd11;
        rom[541][30] = -8'd58;
        rom[541][31] = 8'd31;
        rom[541][32] = 8'd28;
        rom[541][33] = 8'd31;
        rom[541][34] = 8'd38;
        rom[541][35] = -8'd44;
        rom[541][36] = -8'd1;
        rom[541][37] = -8'd22;
        rom[541][38] = -8'd20;
        rom[541][39] = -8'd21;
        rom[541][40] = -8'd26;
        rom[541][41] = 8'd4;
        rom[541][42] = 8'd1;
        rom[541][43] = -8'd38;
        rom[541][44] = 8'd20;
        rom[541][45] = 8'd21;
        rom[541][46] = 8'd10;
        rom[541][47] = -8'd29;
        rom[541][48] = -8'd35;
        rom[541][49] = -8'd2;
        rom[541][50] = 8'd7;
        rom[541][51] = -8'd41;
        rom[541][52] = 8'd31;
        rom[541][53] = 8'd29;
        rom[541][54] = 8'd22;
        rom[541][55] = 8'd70;
        rom[541][56] = -8'd15;
        rom[541][57] = -8'd1;
        rom[541][58] = -8'd41;
        rom[541][59] = -8'd16;
        rom[541][60] = 8'd25;
        rom[541][61] = 8'd18;
        rom[541][62] = -8'd20;
        rom[541][63] = -8'd12;
        rom[542][0] = 8'd32;
        rom[542][1] = -8'd16;
        rom[542][2] = 8'd49;
        rom[542][3] = -8'd19;
        rom[542][4] = -8'd42;
        rom[542][5] = 8'd0;
        rom[542][6] = 8'd7;
        rom[542][7] = 8'd19;
        rom[542][8] = 8'd5;
        rom[542][9] = -8'd29;
        rom[542][10] = -8'd12;
        rom[542][11] = 8'd22;
        rom[542][12] = 8'd14;
        rom[542][13] = -8'd5;
        rom[542][14] = -8'd6;
        rom[542][15] = 8'd23;
        rom[542][16] = -8'd14;
        rom[542][17] = -8'd9;
        rom[542][18] = -8'd20;
        rom[542][19] = -8'd16;
        rom[542][20] = 8'd5;
        rom[542][21] = 8'd24;
        rom[542][22] = 8'd0;
        rom[542][23] = 8'd35;
        rom[542][24] = 8'd11;
        rom[542][25] = 8'd35;
        rom[542][26] = -8'd13;
        rom[542][27] = 8'd17;
        rom[542][28] = -8'd34;
        rom[542][29] = -8'd41;
        rom[542][30] = -8'd1;
        rom[542][31] = -8'd49;
        rom[542][32] = -8'd33;
        rom[542][33] = -8'd10;
        rom[542][34] = -8'd39;
        rom[542][35] = 8'd41;
        rom[542][36] = -8'd58;
        rom[542][37] = -8'd35;
        rom[542][38] = -8'd30;
        rom[542][39] = 8'd19;
        rom[542][40] = 8'd22;
        rom[542][41] = -8'd17;
        rom[542][42] = -8'd5;
        rom[542][43] = 8'd27;
        rom[542][44] = -8'd28;
        rom[542][45] = -8'd31;
        rom[542][46] = 8'd23;
        rom[542][47] = -8'd44;
        rom[542][48] = 8'd26;
        rom[542][49] = -8'd17;
        rom[542][50] = 8'd36;
        rom[542][51] = 8'd33;
        rom[542][52] = 8'd17;
        rom[542][53] = 8'd22;
        rom[542][54] = 8'd1;
        rom[542][55] = 8'd16;
        rom[542][56] = -8'd27;
        rom[542][57] = -8'd45;
        rom[542][58] = 8'd7;
        rom[542][59] = 8'd1;
        rom[542][60] = 8'd15;
        rom[542][61] = 8'd9;
        rom[542][62] = 8'd17;
        rom[542][63] = 8'd24;
        rom[543][0] = -8'd12;
        rom[543][1] = 8'd6;
        rom[543][2] = -8'd40;
        rom[543][3] = 8'd6;
        rom[543][4] = -8'd44;
        rom[543][5] = -8'd5;
        rom[543][6] = -8'd76;
        rom[543][7] = -8'd16;
        rom[543][8] = -8'd5;
        rom[543][9] = 8'd4;
        rom[543][10] = -8'd30;
        rom[543][11] = -8'd27;
        rom[543][12] = -8'd12;
        rom[543][13] = 8'd37;
        rom[543][14] = 8'd2;
        rom[543][15] = 8'd1;
        rom[543][16] = -8'd29;
        rom[543][17] = 8'd23;
        rom[543][18] = -8'd48;
        rom[543][19] = -8'd6;
        rom[543][20] = 8'd0;
        rom[543][21] = 8'd9;
        rom[543][22] = 8'd3;
        rom[543][23] = -8'd2;
        rom[543][24] = 8'd0;
        rom[543][25] = -8'd46;
        rom[543][26] = -8'd11;
        rom[543][27] = 8'd10;
        rom[543][28] = 8'd17;
        rom[543][29] = -8'd9;
        rom[543][30] = 8'd31;
        rom[543][31] = -8'd13;
        rom[543][32] = -8'd22;
        rom[543][33] = -8'd46;
        rom[543][34] = -8'd1;
        rom[543][35] = 8'd8;
        rom[543][36] = -8'd7;
        rom[543][37] = 8'd18;
        rom[543][38] = 8'd3;
        rom[543][39] = -8'd68;
        rom[543][40] = -8'd1;
        rom[543][41] = -8'd5;
        rom[543][42] = -8'd34;
        rom[543][43] = -8'd15;
        rom[543][44] = -8'd8;
        rom[543][45] = -8'd27;
        rom[543][46] = -8'd42;
        rom[543][47] = 8'd8;
        rom[543][48] = -8'd28;
        rom[543][49] = 8'd20;
        rom[543][50] = -8'd22;
        rom[543][51] = -8'd6;
        rom[543][52] = 8'd9;
        rom[543][53] = 8'd4;
        rom[543][54] = -8'd14;
        rom[543][55] = -8'd3;
        rom[543][56] = 8'd6;
        rom[543][57] = -8'd40;
        rom[543][58] = -8'd18;
        rom[543][59] = 8'd20;
        rom[543][60] = -8'd10;
        rom[543][61] = 8'd8;
        rom[543][62] = 8'd3;
        rom[543][63] = -8'd1;
        rom[544][0] = 8'd11;
        rom[544][1] = 8'd1;
        rom[544][2] = 8'd11;
        rom[544][3] = -8'd21;
        rom[544][4] = 8'd10;
        rom[544][5] = 8'd24;
        rom[544][6] = 8'd41;
        rom[544][7] = 8'd12;
        rom[544][8] = -8'd11;
        rom[544][9] = 8'd26;
        rom[544][10] = -8'd41;
        rom[544][11] = 8'd47;
        rom[544][12] = -8'd45;
        rom[544][13] = 8'd4;
        rom[544][14] = 8'd8;
        rom[544][15] = -8'd15;
        rom[544][16] = -8'd7;
        rom[544][17] = -8'd1;
        rom[544][18] = -8'd14;
        rom[544][19] = 8'd14;
        rom[544][20] = -8'd5;
        rom[544][21] = 8'd8;
        rom[544][22] = -8'd67;
        rom[544][23] = -8'd7;
        rom[544][24] = 8'd36;
        rom[544][25] = -8'd17;
        rom[544][26] = 8'd36;
        rom[544][27] = -8'd27;
        rom[544][28] = 8'd10;
        rom[544][29] = 8'd16;
        rom[544][30] = 8'd10;
        rom[544][31] = 8'd18;
        rom[544][32] = -8'd2;
        rom[544][33] = -8'd3;
        rom[544][34] = 8'd21;
        rom[544][35] = 8'd10;
        rom[544][36] = 8'd22;
        rom[544][37] = -8'd5;
        rom[544][38] = -8'd3;
        rom[544][39] = 8'd18;
        rom[544][40] = 8'd13;
        rom[544][41] = 8'd8;
        rom[544][42] = 8'd54;
        rom[544][43] = -8'd46;
        rom[544][44] = -8'd12;
        rom[544][45] = 8'd42;
        rom[544][46] = -8'd36;
        rom[544][47] = 8'd13;
        rom[544][48] = -8'd21;
        rom[544][49] = -8'd63;
        rom[544][50] = 8'd26;
        rom[544][51] = -8'd18;
        rom[544][52] = -8'd20;
        rom[544][53] = 8'd3;
        rom[544][54] = -8'd4;
        rom[544][55] = 8'd18;
        rom[544][56] = -8'd3;
        rom[544][57] = 8'd16;
        rom[544][58] = 8'd26;
        rom[544][59] = 8'd5;
        rom[544][60] = 8'd38;
        rom[544][61] = -8'd13;
        rom[544][62] = 8'd17;
        rom[544][63] = -8'd16;
        rom[545][0] = 8'd0;
        rom[545][1] = -8'd23;
        rom[545][2] = -8'd20;
        rom[545][3] = -8'd58;
        rom[545][4] = -8'd42;
        rom[545][5] = 8'd23;
        rom[545][6] = 8'd60;
        rom[545][7] = 8'd11;
        rom[545][8] = -8'd11;
        rom[545][9] = -8'd53;
        rom[545][10] = 8'd22;
        rom[545][11] = 8'd35;
        rom[545][12] = -8'd17;
        rom[545][13] = 8'd32;
        rom[545][14] = -8'd2;
        rom[545][15] = 8'd19;
        rom[545][16] = 8'd47;
        rom[545][17] = -8'd7;
        rom[545][18] = -8'd15;
        rom[545][19] = 8'd15;
        rom[545][20] = 8'd0;
        rom[545][21] = -8'd8;
        rom[545][22] = -8'd25;
        rom[545][23] = 8'd20;
        rom[545][24] = -8'd21;
        rom[545][25] = -8'd26;
        rom[545][26] = -8'd23;
        rom[545][27] = 8'd7;
        rom[545][28] = 8'd11;
        rom[545][29] = 8'd18;
        rom[545][30] = -8'd18;
        rom[545][31] = -8'd43;
        rom[545][32] = 8'd7;
        rom[545][33] = 8'd37;
        rom[545][34] = 8'd3;
        rom[545][35] = -8'd26;
        rom[545][36] = 8'd6;
        rom[545][37] = -8'd12;
        rom[545][38] = 8'd23;
        rom[545][39] = -8'd47;
        rom[545][40] = 8'd25;
        rom[545][41] = -8'd24;
        rom[545][42] = -8'd38;
        rom[545][43] = 8'd19;
        rom[545][44] = -8'd18;
        rom[545][45] = -8'd13;
        rom[545][46] = -8'd28;
        rom[545][47] = 8'd12;
        rom[545][48] = -8'd46;
        rom[545][49] = -8'd33;
        rom[545][50] = -8'd15;
        rom[545][51] = -8'd60;
        rom[545][52] = -8'd7;
        rom[545][53] = 8'd4;
        rom[545][54] = 8'd37;
        rom[545][55] = 8'd38;
        rom[545][56] = 8'd36;
        rom[545][57] = 8'd6;
        rom[545][58] = 8'd16;
        rom[545][59] = -8'd30;
        rom[545][60] = 8'd23;
        rom[545][61] = -8'd9;
        rom[545][62] = 8'd22;
        rom[545][63] = -8'd7;
        rom[546][0] = 8'd6;
        rom[546][1] = -8'd12;
        rom[546][2] = -8'd47;
        rom[546][3] = -8'd22;
        rom[546][4] = -8'd15;
        rom[546][5] = -8'd3;
        rom[546][6] = -8'd35;
        rom[546][7] = 8'd9;
        rom[546][8] = 8'd42;
        rom[546][9] = -8'd38;
        rom[546][10] = -8'd33;
        rom[546][11] = -8'd27;
        rom[546][12] = -8'd28;
        rom[546][13] = 8'd23;
        rom[546][14] = -8'd10;
        rom[546][15] = -8'd10;
        rom[546][16] = -8'd14;
        rom[546][17] = -8'd17;
        rom[546][18] = 8'd9;
        rom[546][19] = -8'd7;
        rom[546][20] = -8'd2;
        rom[546][21] = 8'd0;
        rom[546][22] = 8'd19;
        rom[546][23] = 8'd19;
        rom[546][24] = 8'd16;
        rom[546][25] = 8'd63;
        rom[546][26] = -8'd2;
        rom[546][27] = 8'd8;
        rom[546][28] = -8'd35;
        rom[546][29] = -8'd3;
        rom[546][30] = 8'd3;
        rom[546][31] = -8'd2;
        rom[546][32] = -8'd39;
        rom[546][33] = 8'd30;
        rom[546][34] = 8'd8;
        rom[546][35] = 8'd6;
        rom[546][36] = 8'd5;
        rom[546][37] = -8'd50;
        rom[546][38] = -8'd39;
        rom[546][39] = 8'd1;
        rom[546][40] = -8'd21;
        rom[546][41] = 8'd34;
        rom[546][42] = -8'd22;
        rom[546][43] = 8'd1;
        rom[546][44] = -8'd18;
        rom[546][45] = 8'd33;
        rom[546][46] = 8'd1;
        rom[546][47] = 8'd20;
        rom[546][48] = -8'd28;
        rom[546][49] = -8'd36;
        rom[546][50] = -8'd1;
        rom[546][51] = 8'd58;
        rom[546][52] = 8'd36;
        rom[546][53] = 8'd8;
        rom[546][54] = 8'd60;
        rom[546][55] = -8'd30;
        rom[546][56] = 8'd30;
        rom[546][57] = 8'd8;
        rom[546][58] = -8'd12;
        rom[546][59] = 8'd2;
        rom[546][60] = -8'd5;
        rom[546][61] = 8'd13;
        rom[546][62] = 8'd36;
        rom[546][63] = -8'd18;
        rom[547][0] = -8'd42;
        rom[547][1] = 8'd30;
        rom[547][2] = -8'd24;
        rom[547][3] = 8'd19;
        rom[547][4] = -8'd7;
        rom[547][5] = 8'd0;
        rom[547][6] = -8'd36;
        rom[547][7] = 8'd7;
        rom[547][8] = 8'd13;
        rom[547][9] = -8'd51;
        rom[547][10] = 8'd9;
        rom[547][11] = 8'd19;
        rom[547][12] = -8'd10;
        rom[547][13] = -8'd13;
        rom[547][14] = 8'd15;
        rom[547][15] = 8'd14;
        rom[547][16] = -8'd12;
        rom[547][17] = 8'd4;
        rom[547][18] = -8'd8;
        rom[547][19] = 8'd15;
        rom[547][20] = 8'd2;
        rom[547][21] = -8'd45;
        rom[547][22] = 8'd5;
        rom[547][23] = -8'd10;
        rom[547][24] = 8'd14;
        rom[547][25] = -8'd25;
        rom[547][26] = -8'd32;
        rom[547][27] = -8'd44;
        rom[547][28] = 8'd22;
        rom[547][29] = 8'd24;
        rom[547][30] = 8'd23;
        rom[547][31] = -8'd6;
        rom[547][32] = 8'd0;
        rom[547][33] = 8'd26;
        rom[547][34] = -8'd27;
        rom[547][35] = -8'd26;
        rom[547][36] = -8'd12;
        rom[547][37] = 8'd2;
        rom[547][38] = -8'd26;
        rom[547][39] = -8'd50;
        rom[547][40] = 8'd8;
        rom[547][41] = 8'd14;
        rom[547][42] = 8'd42;
        rom[547][43] = 8'd20;
        rom[547][44] = 8'd21;
        rom[547][45] = 8'd18;
        rom[547][46] = -8'd56;
        rom[547][47] = -8'd31;
        rom[547][48] = 8'd9;
        rom[547][49] = -8'd14;
        rom[547][50] = 8'd2;
        rom[547][51] = 8'd6;
        rom[547][52] = 8'd12;
        rom[547][53] = -8'd10;
        rom[547][54] = 8'd33;
        rom[547][55] = -8'd23;
        rom[547][56] = 8'd15;
        rom[547][57] = 8'd9;
        rom[547][58] = -8'd18;
        rom[547][59] = -8'd54;
        rom[547][60] = -8'd80;
        rom[547][61] = -8'd21;
        rom[547][62] = -8'd9;
        rom[547][63] = -8'd51;
        rom[548][0] = 8'd12;
        rom[548][1] = -8'd48;
        rom[548][2] = 8'd22;
        rom[548][3] = -8'd3;
        rom[548][4] = -8'd52;
        rom[548][5] = 8'd6;
        rom[548][6] = 8'd50;
        rom[548][7] = -8'd21;
        rom[548][8] = 8'd3;
        rom[548][9] = -8'd34;
        rom[548][10] = -8'd3;
        rom[548][11] = 8'd15;
        rom[548][12] = -8'd35;
        rom[548][13] = -8'd34;
        rom[548][14] = 8'd18;
        rom[548][15] = -8'd26;
        rom[548][16] = -8'd45;
        rom[548][17] = 8'd19;
        rom[548][18] = 8'd14;
        rom[548][19] = -8'd2;
        rom[548][20] = -8'd15;
        rom[548][21] = -8'd13;
        rom[548][22] = -8'd18;
        rom[548][23] = -8'd9;
        rom[548][24] = 8'd1;
        rom[548][25] = -8'd15;
        rom[548][26] = -8'd1;
        rom[548][27] = 8'd27;
        rom[548][28] = 8'd22;
        rom[548][29] = 8'd0;
        rom[548][30] = 8'd6;
        rom[548][31] = 8'd1;
        rom[548][32] = -8'd5;
        rom[548][33] = -8'd7;
        rom[548][34] = -8'd13;
        rom[548][35] = -8'd34;
        rom[548][36] = 8'd10;
        rom[548][37] = -8'd29;
        rom[548][38] = -8'd18;
        rom[548][39] = 8'd16;
        rom[548][40] = 8'd21;
        rom[548][41] = 8'd3;
        rom[548][42] = -8'd3;
        rom[548][43] = -8'd14;
        rom[548][44] = -8'd18;
        rom[548][45] = -8'd37;
        rom[548][46] = -8'd46;
        rom[548][47] = 8'd34;
        rom[548][48] = -8'd19;
        rom[548][49] = 8'd40;
        rom[548][50] = 8'd24;
        rom[548][51] = 8'd17;
        rom[548][52] = -8'd31;
        rom[548][53] = 8'd8;
        rom[548][54] = -8'd7;
        rom[548][55] = -8'd19;
        rom[548][56] = -8'd34;
        rom[548][57] = -8'd3;
        rom[548][58] = 8'd24;
        rom[548][59] = -8'd24;
        rom[548][60] = -8'd41;
        rom[548][61] = -8'd18;
        rom[548][62] = -8'd16;
        rom[548][63] = 8'd2;
        rom[549][0] = 8'd46;
        rom[549][1] = -8'd9;
        rom[549][2] = -8'd47;
        rom[549][3] = 8'd0;
        rom[549][4] = 8'd42;
        rom[549][5] = -8'd12;
        rom[549][6] = -8'd23;
        rom[549][7] = -8'd18;
        rom[549][8] = 8'd5;
        rom[549][9] = 8'd6;
        rom[549][10] = -8'd38;
        rom[549][11] = 8'd38;
        rom[549][12] = 8'd0;
        rom[549][13] = 8'd13;
        rom[549][14] = 8'd16;
        rom[549][15] = -8'd22;
        rom[549][16] = -8'd15;
        rom[549][17] = -8'd38;
        rom[549][18] = 8'd13;
        rom[549][19] = -8'd53;
        rom[549][20] = -8'd7;
        rom[549][21] = -8'd36;
        rom[549][22] = -8'd23;
        rom[549][23] = 8'd55;
        rom[549][24] = 8'd5;
        rom[549][25] = -8'd17;
        rom[549][26] = 8'd14;
        rom[549][27] = -8'd30;
        rom[549][28] = 8'd16;
        rom[549][29] = 8'd15;
        rom[549][30] = -8'd41;
        rom[549][31] = -8'd10;
        rom[549][32] = 8'd22;
        rom[549][33] = -8'd30;
        rom[549][34] = -8'd14;
        rom[549][35] = -8'd66;
        rom[549][36] = -8'd7;
        rom[549][37] = -8'd1;
        rom[549][38] = -8'd12;
        rom[549][39] = -8'd43;
        rom[549][40] = -8'd33;
        rom[549][41] = -8'd9;
        rom[549][42] = -8'd1;
        rom[549][43] = 8'd15;
        rom[549][44] = -8'd3;
        rom[549][45] = 8'd16;
        rom[549][46] = -8'd25;
        rom[549][47] = -8'd19;
        rom[549][48] = -8'd1;
        rom[549][49] = -8'd28;
        rom[549][50] = 8'd24;
        rom[549][51] = -8'd42;
        rom[549][52] = 8'd21;
        rom[549][53] = 8'd31;
        rom[549][54] = -8'd70;
        rom[549][55] = -8'd20;
        rom[549][56] = -8'd45;
        rom[549][57] = -8'd13;
        rom[549][58] = -8'd28;
        rom[549][59] = -8'd20;
        rom[549][60] = -8'd3;
        rom[549][61] = 8'd1;
        rom[549][62] = 8'd24;
        rom[549][63] = 8'd5;
        rom[550][0] = -8'd53;
        rom[550][1] = -8'd40;
        rom[550][2] = -8'd11;
        rom[550][3] = 8'd41;
        rom[550][4] = 8'd12;
        rom[550][5] = -8'd43;
        rom[550][6] = -8'd45;
        rom[550][7] = 8'd16;
        rom[550][8] = 8'd13;
        rom[550][9] = 8'd8;
        rom[550][10] = -8'd29;
        rom[550][11] = 8'd18;
        rom[550][12] = 8'd3;
        rom[550][13] = 8'd3;
        rom[550][14] = -8'd86;
        rom[550][15] = 8'd14;
        rom[550][16] = 8'd30;
        rom[550][17] = -8'd34;
        rom[550][18] = -8'd16;
        rom[550][19] = 8'd2;
        rom[550][20] = -8'd12;
        rom[550][21] = -8'd43;
        rom[550][22] = -8'd13;
        rom[550][23] = 8'd0;
        rom[550][24] = -8'd38;
        rom[550][25] = 8'd17;
        rom[550][26] = -8'd54;
        rom[550][27] = -8'd42;
        rom[550][28] = 8'd51;
        rom[550][29] = 8'd20;
        rom[550][30] = 8'd3;
        rom[550][31] = -8'd12;
        rom[550][32] = 8'd53;
        rom[550][33] = 8'd7;
        rom[550][34] = -8'd25;
        rom[550][35] = -8'd26;
        rom[550][36] = -8'd5;
        rom[550][37] = -8'd74;
        rom[550][38] = -8'd15;
        rom[550][39] = 8'd11;
        rom[550][40] = 8'd30;
        rom[550][41] = 8'd36;
        rom[550][42] = 8'd7;
        rom[550][43] = 8'd6;
        rom[550][44] = 8'd18;
        rom[550][45] = 8'd0;
        rom[550][46] = 8'd2;
        rom[550][47] = -8'd2;
        rom[550][48] = -8'd56;
        rom[550][49] = 8'd13;
        rom[550][50] = 8'd43;
        rom[550][51] = 8'd4;
        rom[550][52] = 8'd23;
        rom[550][53] = -8'd22;
        rom[550][54] = -8'd6;
        rom[550][55] = -8'd35;
        rom[550][56] = 8'd53;
        rom[550][57] = 8'd19;
        rom[550][58] = -8'd16;
        rom[550][59] = 8'd18;
        rom[550][60] = 8'd7;
        rom[550][61] = 8'd14;
        rom[550][62] = -8'd38;
        rom[550][63] = 8'd16;
        rom[551][0] = -8'd8;
        rom[551][1] = -8'd29;
        rom[551][2] = -8'd51;
        rom[551][3] = 8'd47;
        rom[551][4] = 8'd11;
        rom[551][5] = 8'd30;
        rom[551][6] = 8'd3;
        rom[551][7] = 8'd13;
        rom[551][8] = -8'd20;
        rom[551][9] = -8'd2;
        rom[551][10] = -8'd30;
        rom[551][11] = 8'd16;
        rom[551][12] = -8'd27;
        rom[551][13] = 8'd3;
        rom[551][14] = -8'd8;
        rom[551][15] = 8'd34;
        rom[551][16] = -8'd26;
        rom[551][17] = 8'd33;
        rom[551][18] = 8'd9;
        rom[551][19] = -8'd28;
        rom[551][20] = 8'd4;
        rom[551][21] = -8'd29;
        rom[551][22] = -8'd10;
        rom[551][23] = 8'd25;
        rom[551][24] = -8'd30;
        rom[551][25] = -8'd1;
        rom[551][26] = -8'd17;
        rom[551][27] = -8'd68;
        rom[551][28] = -8'd18;
        rom[551][29] = 8'd4;
        rom[551][30] = 8'd36;
        rom[551][31] = 8'd39;
        rom[551][32] = -8'd60;
        rom[551][33] = 8'd6;
        rom[551][34] = -8'd4;
        rom[551][35] = 8'd7;
        rom[551][36] = 8'd15;
        rom[551][37] = -8'd28;
        rom[551][38] = -8'd29;
        rom[551][39] = 8'd14;
        rom[551][40] = -8'd19;
        rom[551][41] = -8'd32;
        rom[551][42] = 8'd4;
        rom[551][43] = 8'd17;
        rom[551][44] = -8'd12;
        rom[551][45] = 8'd18;
        rom[551][46] = -8'd23;
        rom[551][47] = -8'd34;
        rom[551][48] = -8'd44;
        rom[551][49] = 8'd13;
        rom[551][50] = 8'd37;
        rom[551][51] = -8'd22;
        rom[551][52] = 8'd2;
        rom[551][53] = 8'd54;
        rom[551][54] = -8'd17;
        rom[551][55] = -8'd50;
        rom[551][56] = 8'd11;
        rom[551][57] = 8'd38;
        rom[551][58] = -8'd8;
        rom[551][59] = 8'd24;
        rom[551][60] = 8'd5;
        rom[551][61] = 8'd16;
        rom[551][62] = 8'd9;
        rom[551][63] = -8'd6;
        rom[552][0] = 8'd5;
        rom[552][1] = 8'd23;
        rom[552][2] = -8'd21;
        rom[552][3] = -8'd7;
        rom[552][4] = -8'd8;
        rom[552][5] = 8'd1;
        rom[552][6] = 8'd2;
        rom[552][7] = -8'd29;
        rom[552][8] = 8'd30;
        rom[552][9] = 8'd41;
        rom[552][10] = 8'd6;
        rom[552][11] = 8'd18;
        rom[552][12] = -8'd64;
        rom[552][13] = 8'd3;
        rom[552][14] = 8'd26;
        rom[552][15] = -8'd20;
        rom[552][16] = -8'd56;
        rom[552][17] = 8'd23;
        rom[552][18] = 8'd0;
        rom[552][19] = 8'd26;
        rom[552][20] = -8'd11;
        rom[552][21] = 8'd23;
        rom[552][22] = 8'd1;
        rom[552][23] = 8'd18;
        rom[552][24] = -8'd2;
        rom[552][25] = 8'd18;
        rom[552][26] = 8'd6;
        rom[552][27] = -8'd18;
        rom[552][28] = 8'd43;
        rom[552][29] = -8'd20;
        rom[552][30] = 8'd95;
        rom[552][31] = -8'd39;
        rom[552][32] = 8'd22;
        rom[552][33] = -8'd5;
        rom[552][34] = -8'd7;
        rom[552][35] = -8'd1;
        rom[552][36] = 8'd40;
        rom[552][37] = -8'd45;
        rom[552][38] = 8'd1;
        rom[552][39] = 8'd28;
        rom[552][40] = -8'd23;
        rom[552][41] = 8'd33;
        rom[552][42] = -8'd16;
        rom[552][43] = 8'd22;
        rom[552][44] = -8'd18;
        rom[552][45] = 8'd30;
        rom[552][46] = -8'd39;
        rom[552][47] = -8'd1;
        rom[552][48] = -8'd9;
        rom[552][49] = 8'd4;
        rom[552][50] = -8'd42;
        rom[552][51] = 8'd8;
        rom[552][52] = 8'd8;
        rom[552][53] = 8'd4;
        rom[552][54] = -8'd4;
        rom[552][55] = 8'd14;
        rom[552][56] = 8'd25;
        rom[552][57] = 8'd18;
        rom[552][58] = 8'd62;
        rom[552][59] = -8'd22;
        rom[552][60] = 8'd30;
        rom[552][61] = 8'd12;
        rom[552][62] = 8'd23;
        rom[552][63] = 8'd23;
        rom[553][0] = -8'd21;
        rom[553][1] = 8'd14;
        rom[553][2] = -8'd45;
        rom[553][3] = -8'd5;
        rom[553][4] = -8'd66;
        rom[553][5] = -8'd49;
        rom[553][6] = 8'd32;
        rom[553][7] = -8'd89;
        rom[553][8] = 8'd19;
        rom[553][9] = 8'd32;
        rom[553][10] = -8'd25;
        rom[553][11] = -8'd22;
        rom[553][12] = -8'd3;
        rom[553][13] = -8'd8;
        rom[553][14] = 8'd2;
        rom[553][15] = 8'd6;
        rom[553][16] = -8'd78;
        rom[553][17] = -8'd6;
        rom[553][18] = -8'd3;
        rom[553][19] = 8'd15;
        rom[553][20] = -8'd11;
        rom[553][21] = -8'd2;
        rom[553][22] = 8'd31;
        rom[553][23] = -8'd71;
        rom[553][24] = 8'd6;
        rom[553][25] = -8'd3;
        rom[553][26] = -8'd7;
        rom[553][27] = -8'd9;
        rom[553][28] = 8'd2;
        rom[553][29] = -8'd10;
        rom[553][30] = 8'd28;
        rom[553][31] = 8'd37;
        rom[553][32] = 8'd16;
        rom[553][33] = -8'd53;
        rom[553][34] = 8'd40;
        rom[553][35] = -8'd2;
        rom[553][36] = 8'd18;
        rom[553][37] = -8'd21;
        rom[553][38] = -8'd15;
        rom[553][39] = -8'd32;
        rom[553][40] = -8'd54;
        rom[553][41] = 8'd51;
        rom[553][42] = -8'd32;
        rom[553][43] = 8'd15;
        rom[553][44] = -8'd13;
        rom[553][45] = -8'd91;
        rom[553][46] = -8'd14;
        rom[553][47] = -8'd25;
        rom[553][48] = -8'd41;
        rom[553][49] = 8'd68;
        rom[553][50] = 8'd22;
        rom[553][51] = -8'd7;
        rom[553][52] = 8'd6;
        rom[553][53] = 8'd34;
        rom[553][54] = -8'd11;
        rom[553][55] = -8'd13;
        rom[553][56] = -8'd55;
        rom[553][57] = 8'd8;
        rom[553][58] = -8'd25;
        rom[553][59] = -8'd33;
        rom[553][60] = 8'd19;
        rom[553][61] = -8'd64;
        rom[553][62] = -8'd8;
        rom[553][63] = -8'd33;
        rom[554][0] = -8'd25;
        rom[554][1] = -8'd34;
        rom[554][2] = -8'd14;
        rom[554][3] = 8'd36;
        rom[554][4] = 8'd6;
        rom[554][5] = -8'd35;
        rom[554][6] = -8'd14;
        rom[554][7] = 8'd43;
        rom[554][8] = -8'd12;
        rom[554][9] = 8'd9;
        rom[554][10] = -8'd8;
        rom[554][11] = 8'd7;
        rom[554][12] = 8'd7;
        rom[554][13] = 8'd24;
        rom[554][14] = -8'd56;
        rom[554][15] = -8'd17;
        rom[554][16] = 8'd5;
        rom[554][17] = -8'd44;
        rom[554][18] = -8'd1;
        rom[554][19] = -8'd1;
        rom[554][20] = -8'd4;
        rom[554][21] = 8'd14;
        rom[554][22] = 8'd55;
        rom[554][23] = 8'd18;
        rom[554][24] = 8'd26;
        rom[554][25] = -8'd40;
        rom[554][26] = -8'd24;
        rom[554][27] = -8'd63;
        rom[554][28] = 8'd6;
        rom[554][29] = 8'd8;
        rom[554][30] = -8'd35;
        rom[554][31] = 8'd16;
        rom[554][32] = 8'd44;
        rom[554][33] = 8'd41;
        rom[554][34] = -8'd19;
        rom[554][35] = 8'd3;
        rom[554][36] = 8'd0;
        rom[554][37] = 8'd19;
        rom[554][38] = -8'd42;
        rom[554][39] = -8'd13;
        rom[554][40] = -8'd22;
        rom[554][41] = -8'd17;
        rom[554][42] = 8'd20;
        rom[554][43] = 8'd3;
        rom[554][44] = -8'd56;
        rom[554][45] = -8'd37;
        rom[554][46] = 8'd7;
        rom[554][47] = 8'd29;
        rom[554][48] = -8'd1;
        rom[554][49] = 8'd15;
        rom[554][50] = 8'd14;
        rom[554][51] = 8'd40;
        rom[554][52] = -8'd19;
        rom[554][53] = 8'd15;
        rom[554][54] = 8'd10;
        rom[554][55] = 8'd2;
        rom[554][56] = -8'd37;
        rom[554][57] = -8'd58;
        rom[554][58] = 8'd14;
        rom[554][59] = 8'd0;
        rom[554][60] = 8'd31;
        rom[554][61] = 8'd16;
        rom[554][62] = 8'd1;
        rom[554][63] = 8'd2;
        rom[555][0] = -8'd54;
        rom[555][1] = 8'd20;
        rom[555][2] = -8'd49;
        rom[555][3] = -8'd44;
        rom[555][4] = -8'd31;
        rom[555][5] = -8'd6;
        rom[555][6] = 8'd37;
        rom[555][7] = -8'd3;
        rom[555][8] = -8'd13;
        rom[555][9] = 8'd10;
        rom[555][10] = -8'd34;
        rom[555][11] = -8'd5;
        rom[555][12] = -8'd39;
        rom[555][13] = 8'd10;
        rom[555][14] = -8'd14;
        rom[555][15] = -8'd23;
        rom[555][16] = -8'd19;
        rom[555][17] = -8'd15;
        rom[555][18] = -8'd15;
        rom[555][19] = -8'd7;
        rom[555][20] = -8'd4;
        rom[555][21] = -8'd23;
        rom[555][22] = -8'd24;
        rom[555][23] = 8'd1;
        rom[555][24] = -8'd28;
        rom[555][25] = -8'd7;
        rom[555][26] = 8'd4;
        rom[555][27] = -8'd36;
        rom[555][28] = 8'd5;
        rom[555][29] = -8'd5;
        rom[555][30] = 8'd12;
        rom[555][31] = 8'd22;
        rom[555][32] = -8'd2;
        rom[555][33] = -8'd39;
        rom[555][34] = -8'd17;
        rom[555][35] = 8'd9;
        rom[555][36] = -8'd24;
        rom[555][37] = 8'd5;
        rom[555][38] = 8'd61;
        rom[555][39] = 8'd40;
        rom[555][40] = -8'd45;
        rom[555][41] = -8'd41;
        rom[555][42] = -8'd16;
        rom[555][43] = 8'd2;
        rom[555][44] = -8'd8;
        rom[555][45] = 8'd5;
        rom[555][46] = 8'd26;
        rom[555][47] = 8'd33;
        rom[555][48] = -8'd33;
        rom[555][49] = -8'd3;
        rom[555][50] = 8'd15;
        rom[555][51] = -8'd24;
        rom[555][52] = -8'd9;
        rom[555][53] = -8'd14;
        rom[555][54] = 8'd28;
        rom[555][55] = -8'd31;
        rom[555][56] = -8'd23;
        rom[555][57] = -8'd27;
        rom[555][58] = -8'd16;
        rom[555][59] = -8'd18;
        rom[555][60] = -8'd4;
        rom[555][61] = 8'd15;
        rom[555][62] = 8'd6;
        rom[555][63] = 8'd17;
        rom[556][0] = -8'd62;
        rom[556][1] = 8'd14;
        rom[556][2] = -8'd65;
        rom[556][3] = 8'd32;
        rom[556][4] = 8'd9;
        rom[556][5] = 8'd32;
        rom[556][6] = 8'd20;
        rom[556][7] = 8'd7;
        rom[556][8] = -8'd5;
        rom[556][9] = -8'd10;
        rom[556][10] = -8'd48;
        rom[556][11] = 8'd24;
        rom[556][12] = -8'd28;
        rom[556][13] = -8'd41;
        rom[556][14] = -8'd36;
        rom[556][15] = -8'd8;
        rom[556][16] = -8'd11;
        rom[556][17] = 8'd8;
        rom[556][18] = 8'd17;
        rom[556][19] = -8'd19;
        rom[556][20] = 8'd3;
        rom[556][21] = -8'd7;
        rom[556][22] = -8'd46;
        rom[556][23] = -8'd3;
        rom[556][24] = -8'd1;
        rom[556][25] = -8'd18;
        rom[556][26] = -8'd26;
        rom[556][27] = -8'd62;
        rom[556][28] = -8'd12;
        rom[556][29] = -8'd39;
        rom[556][30] = 8'd3;
        rom[556][31] = 8'd58;
        rom[556][32] = -8'd27;
        rom[556][33] = 8'd46;
        rom[556][34] = 8'd40;
        rom[556][35] = 8'd13;
        rom[556][36] = -8'd10;
        rom[556][37] = -8'd3;
        rom[556][38] = 8'd8;
        rom[556][39] = 8'd26;
        rom[556][40] = 8'd58;
        rom[556][41] = -8'd20;
        rom[556][42] = -8'd22;
        rom[556][43] = 8'd15;
        rom[556][44] = 8'd37;
        rom[556][45] = 8'd41;
        rom[556][46] = -8'd42;
        rom[556][47] = -8'd19;
        rom[556][48] = -8'd23;
        rom[556][49] = 8'd31;
        rom[556][50] = 8'd41;
        rom[556][51] = -8'd29;
        rom[556][52] = 8'd10;
        rom[556][53] = 8'd72;
        rom[556][54] = -8'd9;
        rom[556][55] = -8'd15;
        rom[556][56] = -8'd54;
        rom[556][57] = -8'd14;
        rom[556][58] = 8'd3;
        rom[556][59] = -8'd9;
        rom[556][60] = 8'd47;
        rom[556][61] = -8'd12;
        rom[556][62] = -8'd22;
        rom[556][63] = 8'd14;
        rom[557][0] = -8'd23;
        rom[557][1] = 8'd10;
        rom[557][2] = 8'd7;
        rom[557][3] = -8'd21;
        rom[557][4] = 8'd14;
        rom[557][5] = -8'd41;
        rom[557][6] = -8'd88;
        rom[557][7] = 8'd16;
        rom[557][8] = -8'd27;
        rom[557][9] = -8'd63;
        rom[557][10] = 8'd32;
        rom[557][11] = -8'd27;
        rom[557][12] = 8'd31;
        rom[557][13] = -8'd20;
        rom[557][14] = -8'd7;
        rom[557][15] = 8'd12;
        rom[557][16] = -8'd44;
        rom[557][17] = 8'd22;
        rom[557][18] = -8'd12;
        rom[557][19] = 8'd7;
        rom[557][20] = -8'd5;
        rom[557][21] = -8'd21;
        rom[557][22] = 8'd15;
        rom[557][23] = -8'd15;
        rom[557][24] = -8'd22;
        rom[557][25] = -8'd43;
        rom[557][26] = 8'd26;
        rom[557][27] = 8'd42;
        rom[557][28] = 8'd3;
        rom[557][29] = -8'd38;
        rom[557][30] = -8'd28;
        rom[557][31] = -8'd41;
        rom[557][32] = -8'd16;
        rom[557][33] = -8'd57;
        rom[557][34] = -8'd20;
        rom[557][35] = -8'd34;
        rom[557][36] = -8'd16;
        rom[557][37] = -8'd31;
        rom[557][38] = 8'd14;
        rom[557][39] = -8'd29;
        rom[557][40] = -8'd27;
        rom[557][41] = -8'd59;
        rom[557][42] = 8'd40;
        rom[557][43] = -8'd36;
        rom[557][44] = 8'd10;
        rom[557][45] = -8'd69;
        rom[557][46] = -8'd54;
        rom[557][47] = 8'd29;
        rom[557][48] = -8'd24;
        rom[557][49] = 8'd10;
        rom[557][50] = -8'd38;
        rom[557][51] = 8'd32;
        rom[557][52] = -8'd43;
        rom[557][53] = -8'd21;
        rom[557][54] = -8'd20;
        rom[557][55] = 8'd19;
        rom[557][56] = 8'd1;
        rom[557][57] = 8'd1;
        rom[557][58] = -8'd47;
        rom[557][59] = -8'd23;
        rom[557][60] = -8'd10;
        rom[557][61] = 8'd37;
        rom[557][62] = -8'd47;
        rom[557][63] = -8'd4;
        rom[558][0] = 8'd17;
        rom[558][1] = -8'd44;
        rom[558][2] = 8'd9;
        rom[558][3] = 8'd2;
        rom[558][4] = 8'd9;
        rom[558][5] = 8'd4;
        rom[558][6] = 8'd0;
        rom[558][7] = -8'd6;
        rom[558][8] = 8'd0;
        rom[558][9] = -8'd15;
        rom[558][10] = -8'd22;
        rom[558][11] = 8'd20;
        rom[558][12] = -8'd32;
        rom[558][13] = -8'd13;
        rom[558][14] = -8'd6;
        rom[558][15] = 8'd15;
        rom[558][16] = -8'd105;
        rom[558][17] = 8'd8;
        rom[558][18] = 8'd2;
        rom[558][19] = 8'd28;
        rom[558][20] = -8'd3;
        rom[558][21] = -8'd27;
        rom[558][22] = 8'd40;
        rom[558][23] = 8'd25;
        rom[558][24] = 8'd47;
        rom[558][25] = -8'd42;
        rom[558][26] = 8'd21;
        rom[558][27] = -8'd26;
        rom[558][28] = 8'd17;
        rom[558][29] = 8'd3;
        rom[558][30] = -8'd20;
        rom[558][31] = 8'd5;
        rom[558][32] = 8'd5;
        rom[558][33] = -8'd16;
        rom[558][34] = -8'd14;
        rom[558][35] = 8'd12;
        rom[558][36] = 8'd57;
        rom[558][37] = -8'd52;
        rom[558][38] = -8'd5;
        rom[558][39] = -8'd20;
        rom[558][40] = 8'd6;
        rom[558][41] = -8'd6;
        rom[558][42] = -8'd1;
        rom[558][43] = -8'd23;
        rom[558][44] = 8'd14;
        rom[558][45] = -8'd37;
        rom[558][46] = -8'd56;
        rom[558][47] = -8'd30;
        rom[558][48] = 8'd39;
        rom[558][49] = -8'd28;
        rom[558][50] = -8'd75;
        rom[558][51] = 8'd33;
        rom[558][52] = 8'd29;
        rom[558][53] = 8'd10;
        rom[558][54] = 8'd10;
        rom[558][55] = 8'd41;
        rom[558][56] = 8'd17;
        rom[558][57] = -8'd41;
        rom[558][58] = -8'd7;
        rom[558][59] = -8'd51;
        rom[558][60] = 8'd2;
        rom[558][61] = -8'd42;
        rom[558][62] = -8'd29;
        rom[558][63] = -8'd31;
        rom[559][0] = -8'd10;
        rom[559][1] = 8'd49;
        rom[559][2] = -8'd90;
        rom[559][3] = 8'd13;
        rom[559][4] = 8'd19;
        rom[559][5] = 8'd5;
        rom[559][6] = 8'd31;
        rom[559][7] = -8'd22;
        rom[559][8] = -8'd53;
        rom[559][9] = -8'd38;
        rom[559][10] = 8'd6;
        rom[559][11] = -8'd17;
        rom[559][12] = 8'd9;
        rom[559][13] = 8'd67;
        rom[559][14] = 8'd19;
        rom[559][15] = -8'd31;
        rom[559][16] = -8'd15;
        rom[559][17] = 8'd46;
        rom[559][18] = -8'd36;
        rom[559][19] = 8'd18;
        rom[559][20] = -8'd2;
        rom[559][21] = -8'd11;
        rom[559][22] = -8'd17;
        rom[559][23] = -8'd4;
        rom[559][24] = 8'd17;
        rom[559][25] = -8'd9;
        rom[559][26] = -8'd54;
        rom[559][27] = 8'd66;
        rom[559][28] = -8'd24;
        rom[559][29] = -8'd44;
        rom[559][30] = 8'd9;
        rom[559][31] = 8'd6;
        rom[559][32] = -8'd32;
        rom[559][33] = 8'd12;
        rom[559][34] = 8'd53;
        rom[559][35] = 8'd64;
        rom[559][36] = 8'd38;
        rom[559][37] = 8'd33;
        rom[559][38] = 8'd8;
        rom[559][39] = -8'd4;
        rom[559][40] = -8'd20;
        rom[559][41] = -8'd7;
        rom[559][42] = -8'd35;
        rom[559][43] = 8'd13;
        rom[559][44] = 8'd60;
        rom[559][45] = -8'd6;
        rom[559][46] = -8'd58;
        rom[559][47] = 8'd16;
        rom[559][48] = -8'd27;
        rom[559][49] = 8'd25;
        rom[559][50] = -8'd10;
        rom[559][51] = -8'd67;
        rom[559][52] = 8'd0;
        rom[559][53] = -8'd24;
        rom[559][54] = -8'd17;
        rom[559][55] = -8'd33;
        rom[559][56] = -8'd54;
        rom[559][57] = -8'd19;
        rom[559][58] = 8'd42;
        rom[559][59] = -8'd53;
        rom[559][60] = 8'd29;
        rom[559][61] = -8'd5;
        rom[559][62] = -8'd3;
        rom[559][63] = 8'd29;
        rom[560][0] = 8'd3;
        rom[560][1] = -8'd9;
        rom[560][2] = -8'd12;
        rom[560][3] = -8'd6;
        rom[560][4] = 8'd15;
        rom[560][5] = 8'd21;
        rom[560][6] = -8'd25;
        rom[560][7] = 8'd13;
        rom[560][8] = -8'd14;
        rom[560][9] = -8'd17;
        rom[560][10] = -8'd7;
        rom[560][11] = -8'd20;
        rom[560][12] = 8'd49;
        rom[560][13] = 8'd28;
        rom[560][14] = 8'd16;
        rom[560][15] = 8'd22;
        rom[560][16] = -8'd7;
        rom[560][17] = -8'd11;
        rom[560][18] = -8'd43;
        rom[560][19] = 8'd17;
        rom[560][20] = 8'd1;
        rom[560][21] = 8'd0;
        rom[560][22] = 8'd51;
        rom[560][23] = 8'd32;
        rom[560][24] = 8'd2;
        rom[560][25] = 8'd11;
        rom[560][26] = 8'd28;
        rom[560][27] = 8'd20;
        rom[560][28] = -8'd34;
        rom[560][29] = 8'd25;
        rom[560][30] = -8'd50;
        rom[560][31] = -8'd28;
        rom[560][32] = 8'd35;
        rom[560][33] = 8'd13;
        rom[560][34] = 8'd3;
        rom[560][35] = 8'd39;
        rom[560][36] = -8'd15;
        rom[560][37] = -8'd19;
        rom[560][38] = -8'd2;
        rom[560][39] = -8'd34;
        rom[560][40] = 8'd5;
        rom[560][41] = -8'd2;
        rom[560][42] = -8'd31;
        rom[560][43] = -8'd6;
        rom[560][44] = 8'd24;
        rom[560][45] = -8'd39;
        rom[560][46] = 8'd4;
        rom[560][47] = -8'd53;
        rom[560][48] = -8'd44;
        rom[560][49] = 8'd0;
        rom[560][50] = -8'd28;
        rom[560][51] = -8'd99;
        rom[560][52] = -8'd48;
        rom[560][53] = -8'd28;
        rom[560][54] = 8'd3;
        rom[560][55] = -8'd1;
        rom[560][56] = -8'd16;
        rom[560][57] = 8'd5;
        rom[560][58] = 8'd30;
        rom[560][59] = -8'd43;
        rom[560][60] = -8'd1;
        rom[560][61] = 8'd26;
        rom[560][62] = -8'd23;
        rom[560][63] = -8'd4;
        rom[561][0] = -8'd2;
        rom[561][1] = -8'd46;
        rom[561][2] = -8'd60;
        rom[561][3] = 8'd8;
        rom[561][4] = 8'd10;
        rom[561][5] = -8'd17;
        rom[561][6] = 8'd29;
        rom[561][7] = -8'd19;
        rom[561][8] = -8'd27;
        rom[561][9] = -8'd17;
        rom[561][10] = -8'd38;
        rom[561][11] = 8'd32;
        rom[561][12] = 8'd16;
        rom[561][13] = 8'd65;
        rom[561][14] = -8'd20;
        rom[561][15] = -8'd21;
        rom[561][16] = -8'd11;
        rom[561][17] = 8'd4;
        rom[561][18] = 8'd21;
        rom[561][19] = 8'd1;
        rom[561][20] = 8'd2;
        rom[561][21] = -8'd47;
        rom[561][22] = -8'd51;
        rom[561][23] = -8'd3;
        rom[561][24] = 8'd30;
        rom[561][25] = -8'd2;
        rom[561][26] = -8'd13;
        rom[561][27] = 8'd29;
        rom[561][28] = 8'd16;
        rom[561][29] = 8'd15;
        rom[561][30] = -8'd16;
        rom[561][31] = -8'd8;
        rom[561][32] = 8'd12;
        rom[561][33] = 8'd15;
        rom[561][34] = 8'd19;
        rom[561][35] = -8'd1;
        rom[561][36] = 8'd12;
        rom[561][37] = -8'd49;
        rom[561][38] = -8'd24;
        rom[561][39] = -8'd41;
        rom[561][40] = 8'd20;
        rom[561][41] = -8'd46;
        rom[561][42] = -8'd37;
        rom[561][43] = -8'd7;
        rom[561][44] = 8'd25;
        rom[561][45] = 8'd1;
        rom[561][46] = -8'd22;
        rom[561][47] = 8'd5;
        rom[561][48] = -8'd11;
        rom[561][49] = -8'd4;
        rom[561][50] = -8'd15;
        rom[561][51] = -8'd18;
        rom[561][52] = -8'd1;
        rom[561][53] = 8'd15;
        rom[561][54] = -8'd10;
        rom[561][55] = -8'd10;
        rom[561][56] = 8'd19;
        rom[561][57] = -8'd27;
        rom[561][58] = 8'd14;
        rom[561][59] = 8'd14;
        rom[561][60] = -8'd18;
        rom[561][61] = -8'd14;
        rom[561][62] = -8'd35;
        rom[561][63] = 8'd18;
        rom[562][0] = 8'd14;
        rom[562][1] = 8'd5;
        rom[562][2] = 8'd30;
        rom[562][3] = 8'd30;
        rom[562][4] = 8'd23;
        rom[562][5] = -8'd2;
        rom[562][6] = -8'd18;
        rom[562][7] = 8'd1;
        rom[562][8] = 8'd1;
        rom[562][9] = -8'd15;
        rom[562][10] = -8'd25;
        rom[562][11] = 8'd18;
        rom[562][12] = -8'd13;
        rom[562][13] = 8'd24;
        rom[562][14] = -8'd69;
        rom[562][15] = -8'd4;
        rom[562][16] = -8'd37;
        rom[562][17] = -8'd35;
        rom[562][18] = 8'd30;
        rom[562][19] = 8'd8;
        rom[562][20] = -8'd3;
        rom[562][21] = 8'd2;
        rom[562][22] = -8'd2;
        rom[562][23] = -8'd6;
        rom[562][24] = 8'd43;
        rom[562][25] = -8'd31;
        rom[562][26] = -8'd16;
        rom[562][27] = -8'd13;
        rom[562][28] = -8'd24;
        rom[562][29] = -8'd27;
        rom[562][30] = 8'd25;
        rom[562][31] = 8'd7;
        rom[562][32] = 8'd34;
        rom[562][33] = -8'd26;
        rom[562][34] = -8'd24;
        rom[562][35] = 8'd21;
        rom[562][36] = 8'd12;
        rom[562][37] = -8'd73;
        rom[562][38] = 8'd25;
        rom[562][39] = 8'd1;
        rom[562][40] = -8'd9;
        rom[562][41] = 8'd26;
        rom[562][42] = -8'd57;
        rom[562][43] = -8'd30;
        rom[562][44] = -8'd19;
        rom[562][45] = -8'd24;
        rom[562][46] = 8'd21;
        rom[562][47] = 8'd67;
        rom[562][48] = -8'd9;
        rom[562][49] = 8'd26;
        rom[562][50] = 8'd22;
        rom[562][51] = -8'd35;
        rom[562][52] = -8'd54;
        rom[562][53] = -8'd2;
        rom[562][54] = -8'd5;
        rom[562][55] = 8'd37;
        rom[562][56] = 8'd4;
        rom[562][57] = -8'd37;
        rom[562][58] = -8'd39;
        rom[562][59] = -8'd37;
        rom[562][60] = 8'd6;
        rom[562][61] = 8'd41;
        rom[562][62] = 8'd9;
        rom[562][63] = -8'd17;
        rom[563][0] = -8'd18;
        rom[563][1] = -8'd37;
        rom[563][2] = 8'd11;
        rom[563][3] = -8'd4;
        rom[563][4] = -8'd43;
        rom[563][5] = -8'd11;
        rom[563][6] = 8'd0;
        rom[563][7] = -8'd6;
        rom[563][8] = 8'd6;
        rom[563][9] = -8'd24;
        rom[563][10] = -8'd1;
        rom[563][11] = 8'd48;
        rom[563][12] = 8'd14;
        rom[563][13] = -8'd3;
        rom[563][14] = 8'd5;
        rom[563][15] = -8'd48;
        rom[563][16] = 8'd23;
        rom[563][17] = -8'd17;
        rom[563][18] = -8'd24;
        rom[563][19] = -8'd35;
        rom[563][20] = -8'd4;
        rom[563][21] = 8'd24;
        rom[563][22] = 8'd17;
        rom[563][23] = -8'd69;
        rom[563][24] = 8'd5;
        rom[563][25] = -8'd4;
        rom[563][26] = -8'd36;
        rom[563][27] = 8'd13;
        rom[563][28] = -8'd3;
        rom[563][29] = -8'd2;
        rom[563][30] = -8'd9;
        rom[563][31] = -8'd30;
        rom[563][32] = -8'd37;
        rom[563][33] = -8'd45;
        rom[563][34] = 8'd7;
        rom[563][35] = -8'd64;
        rom[563][36] = 8'd15;
        rom[563][37] = -8'd5;
        rom[563][38] = 8'd9;
        rom[563][39] = -8'd34;
        rom[563][40] = -8'd36;
        rom[563][41] = -8'd23;
        rom[563][42] = 8'd14;
        rom[563][43] = -8'd18;
        rom[563][44] = 8'd1;
        rom[563][45] = 8'd18;
        rom[563][46] = -8'd52;
        rom[563][47] = 8'd70;
        rom[563][48] = -8'd26;
        rom[563][49] = -8'd46;
        rom[563][50] = -8'd43;
        rom[563][51] = -8'd12;
        rom[563][52] = 8'd4;
        rom[563][53] = -8'd33;
        rom[563][54] = 8'd48;
        rom[563][55] = 8'd43;
        rom[563][56] = -8'd8;
        rom[563][57] = -8'd47;
        rom[563][58] = 8'd3;
        rom[563][59] = -8'd5;
        rom[563][60] = 8'd13;
        rom[563][61] = 8'd15;
        rom[563][62] = -8'd19;
        rom[563][63] = 8'd13;
        rom[564][0] = 8'd18;
        rom[564][1] = -8'd1;
        rom[564][2] = -8'd13;
        rom[564][3] = -8'd62;
        rom[564][4] = -8'd4;
        rom[564][5] = 8'd37;
        rom[564][6] = -8'd31;
        rom[564][7] = 8'd22;
        rom[564][8] = -8'd33;
        rom[564][9] = 8'd13;
        rom[564][10] = -8'd22;
        rom[564][11] = 8'd24;
        rom[564][12] = -8'd36;
        rom[564][13] = 8'd44;
        rom[564][14] = -8'd22;
        rom[564][15] = -8'd12;
        rom[564][16] = -8'd10;
        rom[564][17] = -8'd20;
        rom[564][18] = 8'd11;
        rom[564][19] = -8'd9;
        rom[564][20] = -8'd1;
        rom[564][21] = 8'd37;
        rom[564][22] = -8'd92;
        rom[564][23] = 8'd30;
        rom[564][24] = 8'd7;
        rom[564][25] = -8'd41;
        rom[564][26] = 8'd12;
        rom[564][27] = 8'd42;
        rom[564][28] = 8'd44;
        rom[564][29] = 8'd5;
        rom[564][30] = 8'd18;
        rom[564][31] = -8'd11;
        rom[564][32] = 8'd24;
        rom[564][33] = 8'd36;
        rom[564][34] = -8'd11;
        rom[564][35] = -8'd29;
        rom[564][36] = 8'd37;
        rom[564][37] = 8'd59;
        rom[564][38] = -8'd20;
        rom[564][39] = 8'd46;
        rom[564][40] = 8'd31;
        rom[564][41] = -8'd26;
        rom[564][42] = -8'd43;
        rom[564][43] = -8'd53;
        rom[564][44] = 8'd25;
        rom[564][45] = -8'd2;
        rom[564][46] = -8'd12;
        rom[564][47] = -8'd11;
        rom[564][48] = -8'd18;
        rom[564][49] = 8'd9;
        rom[564][50] = 8'd24;
        rom[564][51] = -8'd65;
        rom[564][52] = 8'd39;
        rom[564][53] = 8'd14;
        rom[564][54] = -8'd51;
        rom[564][55] = 8'd16;
        rom[564][56] = 8'd14;
        rom[564][57] = -8'd30;
        rom[564][58] = 8'd19;
        rom[564][59] = -8'd34;
        rom[564][60] = -8'd45;
        rom[564][61] = -8'd6;
        rom[564][62] = 8'd37;
        rom[564][63] = -8'd32;
        rom[565][0] = 8'd3;
        rom[565][1] = -8'd17;
        rom[565][2] = 8'd1;
        rom[565][3] = -8'd37;
        rom[565][4] = 8'd25;
        rom[565][5] = -8'd29;
        rom[565][6] = -8'd1;
        rom[565][7] = 8'd51;
        rom[565][8] = 8'd3;
        rom[565][9] = 8'd0;
        rom[565][10] = 8'd9;
        rom[565][11] = -8'd32;
        rom[565][12] = -8'd15;
        rom[565][13] = 8'd2;
        rom[565][14] = 8'd41;
        rom[565][15] = -8'd14;
        rom[565][16] = 8'd17;
        rom[565][17] = -8'd69;
        rom[565][18] = -8'd23;
        rom[565][19] = -8'd85;
        rom[565][20] = 8'd0;
        rom[565][21] = 8'd22;
        rom[565][22] = 8'd41;
        rom[565][23] = -8'd17;
        rom[565][24] = 8'd12;
        rom[565][25] = -8'd12;
        rom[565][26] = -8'd23;
        rom[565][27] = 8'd2;
        rom[565][28] = 8'd5;
        rom[565][29] = -8'd18;
        rom[565][30] = -8'd15;
        rom[565][31] = -8'd27;
        rom[565][32] = 8'd45;
        rom[565][33] = -8'd27;
        rom[565][34] = -8'd14;
        rom[565][35] = -8'd23;
        rom[565][36] = -8'd47;
        rom[565][37] = -8'd1;
        rom[565][38] = -8'd28;
        rom[565][39] = 8'd7;
        rom[565][40] = 8'd19;
        rom[565][41] = 8'd6;
        rom[565][42] = -8'd18;
        rom[565][43] = 8'd29;
        rom[565][44] = 8'd11;
        rom[565][45] = -8'd38;
        rom[565][46] = -8'd5;
        rom[565][47] = -8'd21;
        rom[565][48] = 8'd10;
        rom[565][49] = 8'd33;
        rom[565][50] = -8'd33;
        rom[565][51] = 8'd16;
        rom[565][52] = 8'd38;
        rom[565][53] = 8'd14;
        rom[565][54] = 8'd29;
        rom[565][55] = -8'd11;
        rom[565][56] = 8'd12;
        rom[565][57] = -8'd30;
        rom[565][58] = -8'd12;
        rom[565][59] = -8'd16;
        rom[565][60] = 8'd27;
        rom[565][61] = 8'd15;
        rom[565][62] = -8'd33;
        rom[565][63] = -8'd24;
        rom[566][0] = -8'd9;
        rom[566][1] = 8'd1;
        rom[566][2] = -8'd1;
        rom[566][3] = -8'd5;
        rom[566][4] = 8'd6;
        rom[566][5] = 8'd5;
        rom[566][6] = -8'd8;
        rom[566][7] = -8'd7;
        rom[566][8] = -8'd3;
        rom[566][9] = 8'd3;
        rom[566][10] = -8'd8;
        rom[566][11] = -8'd8;
        rom[566][12] = 8'd4;
        rom[566][13] = 8'd4;
        rom[566][14] = -8'd5;
        rom[566][15] = -8'd8;
        rom[566][16] = -8'd9;
        rom[566][17] = 8'd4;
        rom[566][18] = -8'd11;
        rom[566][19] = -8'd1;
        rom[566][20] = -8'd5;
        rom[566][21] = -8'd13;
        rom[566][22] = -8'd1;
        rom[566][23] = -8'd3;
        rom[566][24] = -8'd8;
        rom[566][25] = -8'd2;
        rom[566][26] = 8'd0;
        rom[566][27] = 8'd6;
        rom[566][28] = 8'd0;
        rom[566][29] = 8'd4;
        rom[566][30] = -8'd15;
        rom[566][31] = 8'd1;
        rom[566][32] = -8'd9;
        rom[566][33] = 8'd1;
        rom[566][34] = -8'd8;
        rom[566][35] = 8'd1;
        rom[566][36] = -8'd9;
        rom[566][37] = 8'd0;
        rom[566][38] = 8'd4;
        rom[566][39] = 8'd6;
        rom[566][40] = -8'd6;
        rom[566][41] = -8'd4;
        rom[566][42] = 8'd8;
        rom[566][43] = -8'd6;
        rom[566][44] = -8'd10;
        rom[566][45] = -8'd2;
        rom[566][46] = 8'd2;
        rom[566][47] = 8'd13;
        rom[566][48] = 8'd5;
        rom[566][49] = 8'd6;
        rom[566][50] = -8'd7;
        rom[566][51] = -8'd4;
        rom[566][52] = 8'd2;
        rom[566][53] = 8'd15;
        rom[566][54] = -8'd11;
        rom[566][55] = -8'd13;
        rom[566][56] = 8'd3;
        rom[566][57] = -8'd4;
        rom[566][58] = -8'd2;
        rom[566][59] = 8'd8;
        rom[566][60] = 8'd9;
        rom[566][61] = 8'd2;
        rom[566][62] = 8'd6;
        rom[566][63] = -8'd1;
        rom[567][0] = -8'd69;
        rom[567][1] = -8'd7;
        rom[567][2] = -8'd78;
        rom[567][3] = -8'd6;
        rom[567][4] = -8'd40;
        rom[567][5] = 8'd17;
        rom[567][6] = -8'd65;
        rom[567][7] = 8'd21;
        rom[567][8] = -8'd56;
        rom[567][9] = -8'd26;
        rom[567][10] = -8'd57;
        rom[567][11] = -8'd23;
        rom[567][12] = 8'd5;
        rom[567][13] = 8'd6;
        rom[567][14] = -8'd42;
        rom[567][15] = -8'd29;
        rom[567][16] = -8'd5;
        rom[567][17] = -8'd31;
        rom[567][18] = -8'd14;
        rom[567][19] = -8'd54;
        rom[567][20] = -8'd10;
        rom[567][21] = -8'd25;
        rom[567][22] = -8'd67;
        rom[567][23] = -8'd29;
        rom[567][24] = 8'd13;
        rom[567][25] = -8'd28;
        rom[567][26] = 8'd8;
        rom[567][27] = 8'd7;
        rom[567][28] = -8'd35;
        rom[567][29] = 8'd53;
        rom[567][30] = 8'd1;
        rom[567][31] = -8'd15;
        rom[567][32] = -8'd47;
        rom[567][33] = 8'd13;
        rom[567][34] = -8'd2;
        rom[567][35] = -8'd14;
        rom[567][36] = -8'd26;
        rom[567][37] = -8'd1;
        rom[567][38] = -8'd29;
        rom[567][39] = 8'd17;
        rom[567][40] = 8'd42;
        rom[567][41] = -8'd11;
        rom[567][42] = 8'd8;
        rom[567][43] = 8'd0;
        rom[567][44] = 8'd11;
        rom[567][45] = -8'd12;
        rom[567][46] = -8'd23;
        rom[567][47] = 8'd19;
        rom[567][48] = -8'd47;
        rom[567][49] = 8'd6;
        rom[567][50] = 8'd10;
        rom[567][51] = -8'd7;
        rom[567][52] = -8'd2;
        rom[567][53] = 8'd36;
        rom[567][54] = -8'd35;
        rom[567][55] = -8'd46;
        rom[567][56] = -8'd13;
        rom[567][57] = 8'd18;
        rom[567][58] = -8'd17;
        rom[567][59] = 8'd20;
        rom[567][60] = -8'd24;
        rom[567][61] = 8'd9;
        rom[567][62] = 8'd5;
        rom[567][63] = -8'd34;
        rom[568][0] = -8'd57;
        rom[568][1] = -8'd28;
        rom[568][2] = 8'd10;
        rom[568][3] = 8'd22;
        rom[568][4] = 8'd14;
        rom[568][5] = -8'd15;
        rom[568][6] = -8'd52;
        rom[568][7] = -8'd9;
        rom[568][8] = 8'd10;
        rom[568][9] = 8'd19;
        rom[568][10] = -8'd36;
        rom[568][11] = -8'd22;
        rom[568][12] = 8'd31;
        rom[568][13] = -8'd7;
        rom[568][14] = -8'd67;
        rom[568][15] = -8'd36;
        rom[568][16] = -8'd3;
        rom[568][17] = -8'd16;
        rom[568][18] = -8'd53;
        rom[568][19] = -8'd8;
        rom[568][20] = 8'd4;
        rom[568][21] = 8'd1;
        rom[568][22] = -8'd17;
        rom[568][23] = 8'd1;
        rom[568][24] = 8'd46;
        rom[568][25] = -8'd45;
        rom[568][26] = -8'd72;
        rom[568][27] = 8'd29;
        rom[568][28] = 8'd33;
        rom[568][29] = -8'd11;
        rom[568][30] = 8'd23;
        rom[568][31] = -8'd93;
        rom[568][32] = -8'd8;
        rom[568][33] = -8'd28;
        rom[568][34] = -8'd11;
        rom[568][35] = 8'd14;
        rom[568][36] = -8'd8;
        rom[568][37] = -8'd21;
        rom[568][38] = 8'd25;
        rom[568][39] = -8'd8;
        rom[568][40] = 8'd28;
        rom[568][41] = 8'd45;
        rom[568][42] = -8'd21;
        rom[568][43] = -8'd29;
        rom[568][44] = -8'd19;
        rom[568][45] = 8'd10;
        rom[568][46] = -8'd5;
        rom[568][47] = 8'd8;
        rom[568][48] = -8'd35;
        rom[568][49] = -8'd5;
        rom[568][50] = -8'd16;
        rom[568][51] = -8'd30;
        rom[568][52] = 8'd11;
        rom[568][53] = 8'd13;
        rom[568][54] = 8'd26;
        rom[568][55] = 8'd28;
        rom[568][56] = -8'd41;
        rom[568][57] = 8'd4;
        rom[568][58] = -8'd10;
        rom[568][59] = 8'd1;
        rom[568][60] = -8'd17;
        rom[568][61] = 8'd5;
        rom[568][62] = 8'd15;
        rom[568][63] = 8'd13;
        rom[569][0] = -8'd8;
        rom[569][1] = 8'd34;
        rom[569][2] = -8'd23;
        rom[569][3] = -8'd2;
        rom[569][4] = 8'd38;
        rom[569][5] = 8'd10;
        rom[569][6] = -8'd29;
        rom[569][7] = 8'd27;
        rom[569][8] = -8'd49;
        rom[569][9] = 8'd47;
        rom[569][10] = -8'd34;
        rom[569][11] = 8'd27;
        rom[569][12] = 8'd20;
        rom[569][13] = -8'd5;
        rom[569][14] = -8'd20;
        rom[569][15] = 8'd24;
        rom[569][16] = -8'd2;
        rom[569][17] = 8'd15;
        rom[569][18] = 8'd4;
        rom[569][19] = -8'd16;
        rom[569][20] = 8'd3;
        rom[569][21] = -8'd50;
        rom[569][22] = -8'd32;
        rom[569][23] = 8'd2;
        rom[569][24] = 8'd42;
        rom[569][25] = 8'd13;
        rom[569][26] = 8'd18;
        rom[569][27] = -8'd22;
        rom[569][28] = -8'd6;
        rom[569][29] = -8'd21;
        rom[569][30] = 8'd7;
        rom[569][31] = 8'd16;
        rom[569][32] = -8'd26;
        rom[569][33] = 8'd0;
        rom[569][34] = 8'd25;
        rom[569][35] = 8'd28;
        rom[569][36] = -8'd23;
        rom[569][37] = -8'd11;
        rom[569][38] = -8'd20;
        rom[569][39] = -8'd20;
        rom[569][40] = -8'd26;
        rom[569][41] = 8'd7;
        rom[569][42] = 8'd19;
        rom[569][43] = -8'd27;
        rom[569][44] = 8'd18;
        rom[569][45] = -8'd10;
        rom[569][46] = -8'd23;
        rom[569][47] = -8'd54;
        rom[569][48] = 8'd3;
        rom[569][49] = 8'd29;
        rom[569][50] = 8'd10;
        rom[569][51] = -8'd43;
        rom[569][52] = 8'd2;
        rom[569][53] = -8'd29;
        rom[569][54] = 8'd34;
        rom[569][55] = 8'd7;
        rom[569][56] = 8'd10;
        rom[569][57] = -8'd72;
        rom[569][58] = 8'd1;
        rom[569][59] = -8'd6;
        rom[569][60] = -8'd18;
        rom[569][61] = 8'd27;
        rom[569][62] = -8'd63;
        rom[569][63] = 8'd6;
        rom[570][0] = -8'd3;
        rom[570][1] = 8'd33;
        rom[570][2] = 8'd19;
        rom[570][3] = -8'd14;
        rom[570][4] = -8'd29;
        rom[570][5] = -8'd32;
        rom[570][6] = -8'd17;
        rom[570][7] = -8'd4;
        rom[570][8] = -8'd29;
        rom[570][9] = -8'd24;
        rom[570][10] = 8'd38;
        rom[570][11] = -8'd15;
        rom[570][12] = -8'd45;
        rom[570][13] = -8'd28;
        rom[570][14] = 8'd5;
        rom[570][15] = 8'd50;
        rom[570][16] = -8'd50;
        rom[570][17] = 8'd7;
        rom[570][18] = 8'd23;
        rom[570][19] = 8'd6;
        rom[570][20] = 8'd2;
        rom[570][21] = 8'd45;
        rom[570][22] = 8'd4;
        rom[570][23] = -8'd72;
        rom[570][24] = 8'd27;
        rom[570][25] = 8'd0;
        rom[570][26] = 8'd8;
        rom[570][27] = 8'd23;
        rom[570][28] = 8'd11;
        rom[570][29] = -8'd18;
        rom[570][30] = 8'd23;
        rom[570][31] = -8'd14;
        rom[570][32] = -8'd4;
        rom[570][33] = -8'd11;
        rom[570][34] = 8'd11;
        rom[570][35] = -8'd62;
        rom[570][36] = -8'd10;
        rom[570][37] = 8'd4;
        rom[570][38] = -8'd35;
        rom[570][39] = -8'd2;
        rom[570][40] = -8'd39;
        rom[570][41] = 8'd13;
        rom[570][42] = -8'd66;
        rom[570][43] = 8'd25;
        rom[570][44] = -8'd11;
        rom[570][45] = -8'd71;
        rom[570][46] = 8'd16;
        rom[570][47] = -8'd6;
        rom[570][48] = 8'd41;
        rom[570][49] = 8'd59;
        rom[570][50] = -8'd13;
        rom[570][51] = 8'd63;
        rom[570][52] = 8'd16;
        rom[570][53] = 8'd55;
        rom[570][54] = 8'd28;
        rom[570][55] = -8'd16;
        rom[570][56] = 8'd22;
        rom[570][57] = -8'd75;
        rom[570][58] = 8'd0;
        rom[570][59] = -8'd30;
        rom[570][60] = 8'd30;
        rom[570][61] = 8'd15;
        rom[570][62] = -8'd29;
        rom[570][63] = 8'd6;
        rom[571][0] = -8'd33;
        rom[571][1] = 8'd3;
        rom[571][2] = -8'd40;
        rom[571][3] = -8'd33;
        rom[571][4] = -8'd26;
        rom[571][5] = -8'd24;
        rom[571][6] = -8'd24;
        rom[571][7] = -8'd1;
        rom[571][8] = -8'd33;
        rom[571][9] = 8'd4;
        rom[571][10] = -8'd29;
        rom[571][11] = 8'd22;
        rom[571][12] = 8'd28;
        rom[571][13] = 8'd6;
        rom[571][14] = -8'd5;
        rom[571][15] = 8'd2;
        rom[571][16] = 8'd17;
        rom[571][17] = 8'd23;
        rom[571][18] = -8'd19;
        rom[571][19] = -8'd29;
        rom[571][20] = 8'd8;
        rom[571][21] = -8'd36;
        rom[571][22] = -8'd62;
        rom[571][23] = -8'd5;
        rom[571][24] = -8'd6;
        rom[571][25] = -8'd25;
        rom[571][26] = 8'd24;
        rom[571][27] = 8'd3;
        rom[571][28] = 8'd18;
        rom[571][29] = 8'd25;
        rom[571][30] = 8'd29;
        rom[571][31] = 8'd17;
        rom[571][32] = 8'd47;
        rom[571][33] = 8'd9;
        rom[571][34] = -8'd30;
        rom[571][35] = -8'd49;
        rom[571][36] = 8'd14;
        rom[571][37] = -8'd33;
        rom[571][38] = -8'd32;
        rom[571][39] = -8'd21;
        rom[571][40] = 8'd33;
        rom[571][41] = -8'd13;
        rom[571][42] = 8'd10;
        rom[571][43] = -8'd57;
        rom[571][44] = -8'd43;
        rom[571][45] = 8'd42;
        rom[571][46] = 8'd19;
        rom[571][47] = -8'd18;
        rom[571][48] = -8'd20;
        rom[571][49] = 8'd15;
        rom[571][50] = 8'd28;
        rom[571][51] = -8'd29;
        rom[571][52] = -8'd32;
        rom[571][53] = -8'd37;
        rom[571][54] = -8'd10;
        rom[571][55] = -8'd39;
        rom[571][56] = 8'd3;
        rom[571][57] = -8'd8;
        rom[571][58] = -8'd34;
        rom[571][59] = -8'd14;
        rom[571][60] = -8'd47;
        rom[571][61] = 8'd9;
        rom[571][62] = 8'd24;
        rom[571][63] = 8'd24;
        rom[572][0] = 8'd33;
        rom[572][1] = 8'd10;
        rom[572][2] = -8'd11;
        rom[572][3] = -8'd13;
        rom[572][4] = 8'd19;
        rom[572][5] = -8'd46;
        rom[572][6] = -8'd39;
        rom[572][7] = -8'd9;
        rom[572][8] = 8'd2;
        rom[572][9] = -8'd48;
        rom[572][10] = 8'd24;
        rom[572][11] = 8'd14;
        rom[572][12] = -8'd70;
        rom[572][13] = -8'd44;
        rom[572][14] = 8'd12;
        rom[572][15] = 8'd32;
        rom[572][16] = -8'd3;
        rom[572][17] = 8'd21;
        rom[572][18] = -8'd22;
        rom[572][19] = 8'd26;
        rom[572][20] = 8'd0;
        rom[572][21] = -8'd1;
        rom[572][22] = -8'd20;
        rom[572][23] = -8'd21;
        rom[572][24] = 8'd11;
        rom[572][25] = 8'd7;
        rom[572][26] = -8'd38;
        rom[572][27] = 8'd18;
        rom[572][28] = -8'd15;
        rom[572][29] = -8'd18;
        rom[572][30] = 8'd19;
        rom[572][31] = -8'd45;
        rom[572][32] = 8'd37;
        rom[572][33] = 8'd16;
        rom[572][34] = 8'd27;
        rom[572][35] = -8'd22;
        rom[572][36] = 8'd12;
        rom[572][37] = 8'd0;
        rom[572][38] = -8'd33;
        rom[572][39] = 8'd25;
        rom[572][40] = 8'd22;
        rom[572][41] = -8'd9;
        rom[572][42] = 8'd4;
        rom[572][43] = 8'd24;
        rom[572][44] = -8'd17;
        rom[572][45] = 8'd37;
        rom[572][46] = -8'd16;
        rom[572][47] = 8'd20;
        rom[572][48] = 8'd13;
        rom[572][49] = -8'd27;
        rom[572][50] = 8'd57;
        rom[572][51] = -8'd42;
        rom[572][52] = -8'd54;
        rom[572][53] = -8'd40;
        rom[572][54] = -8'd2;
        rom[572][55] = 8'd13;
        rom[572][56] = 8'd13;
        rom[572][57] = -8'd30;
        rom[572][58] = 8'd6;
        rom[572][59] = -8'd49;
        rom[572][60] = 8'd21;
        rom[572][61] = 8'd1;
        rom[572][62] = -8'd5;
        rom[572][63] = 8'd13;
        rom[573][0] = 8'd20;
        rom[573][1] = -8'd14;
        rom[573][2] = 8'd6;
        rom[573][3] = -8'd57;
        rom[573][4] = -8'd8;
        rom[573][5] = -8'd3;
        rom[573][6] = -8'd48;
        rom[573][7] = 8'd7;
        rom[573][8] = -8'd75;
        rom[573][9] = 8'd45;
        rom[573][10] = -8'd22;
        rom[573][11] = -8'd19;
        rom[573][12] = 8'd37;
        rom[573][13] = 8'd28;
        rom[573][14] = -8'd32;
        rom[573][15] = -8'd22;
        rom[573][16] = -8'd14;
        rom[573][17] = -8'd30;
        rom[573][18] = 8'd64;
        rom[573][19] = 8'd12;
        rom[573][20] = -8'd10;
        rom[573][21] = -8'd46;
        rom[573][22] = 8'd9;
        rom[573][23] = 8'd17;
        rom[573][24] = 8'd31;
        rom[573][25] = -8'd46;
        rom[573][26] = -8'd25;
        rom[573][27] = -8'd23;
        rom[573][28] = 8'd1;
        rom[573][29] = -8'd4;
        rom[573][30] = -8'd25;
        rom[573][31] = -8'd16;
        rom[573][32] = 8'd3;
        rom[573][33] = 8'd2;
        rom[573][34] = 8'd37;
        rom[573][35] = 8'd8;
        rom[573][36] = -8'd26;
        rom[573][37] = -8'd48;
        rom[573][38] = -8'd1;
        rom[573][39] = -8'd3;
        rom[573][40] = 8'd26;
        rom[573][41] = 8'd26;
        rom[573][42] = -8'd24;
        rom[573][43] = -8'd2;
        rom[573][44] = 8'd35;
        rom[573][45] = -8'd11;
        rom[573][46] = -8'd11;
        rom[573][47] = 8'd8;
        rom[573][48] = -8'd27;
        rom[573][49] = 8'd27;
        rom[573][50] = -8'd16;
        rom[573][51] = 8'd25;
        rom[573][52] = 8'd6;
        rom[573][53] = 8'd1;
        rom[573][54] = 8'd15;
        rom[573][55] = -8'd8;
        rom[573][56] = -8'd30;
        rom[573][57] = 8'd28;
        rom[573][58] = -8'd42;
        rom[573][59] = 8'd27;
        rom[573][60] = -8'd3;
        rom[573][61] = 8'd1;
        rom[573][62] = -8'd13;
        rom[573][63] = -8'd2;
        rom[574][0] = 8'd13;
        rom[574][1] = -8'd1;
        rom[574][2] = -8'd2;
        rom[574][3] = -8'd17;
        rom[574][4] = -8'd37;
        rom[574][5] = -8'd10;
        rom[574][6] = -8'd13;
        rom[574][7] = 8'd4;
        rom[574][8] = -8'd7;
        rom[574][9] = -8'd11;
        rom[574][10] = -8'd62;
        rom[574][11] = 8'd5;
        rom[574][12] = 8'd21;
        rom[574][13] = 8'd7;
        rom[574][14] = 8'd36;
        rom[574][15] = 8'd1;
        rom[574][16] = 8'd30;
        rom[574][17] = -8'd17;
        rom[574][18] = 8'd25;
        rom[574][19] = 8'd5;
        rom[574][20] = -8'd10;
        rom[574][21] = -8'd12;
        rom[574][22] = -8'd14;
        rom[574][23] = 8'd8;
        rom[574][24] = -8'd8;
        rom[574][25] = -8'd13;
        rom[574][26] = -8'd3;
        rom[574][27] = 8'd13;
        rom[574][28] = -8'd44;
        rom[574][29] = -8'd15;
        rom[574][30] = -8'd37;
        rom[574][31] = -8'd19;
        rom[574][32] = 8'd5;
        rom[574][33] = 8'd32;
        rom[574][34] = 8'd5;
        rom[574][35] = -8'd51;
        rom[574][36] = 8'd9;
        rom[574][37] = -8'd94;
        rom[574][38] = -8'd18;
        rom[574][39] = 8'd18;
        rom[574][40] = -8'd31;
        rom[574][41] = -8'd15;
        rom[574][42] = 8'd36;
        rom[574][43] = 8'd5;
        rom[574][44] = -8'd23;
        rom[574][45] = 8'd8;
        rom[574][46] = 8'd30;
        rom[574][47] = -8'd47;
        rom[574][48] = 8'd8;
        rom[574][49] = -8'd86;
        rom[574][50] = 8'd17;
        rom[574][51] = -8'd43;
        rom[574][52] = 8'd19;
        rom[574][53] = -8'd21;
        rom[574][54] = 8'd27;
        rom[574][55] = -8'd34;
        rom[574][56] = -8'd30;
        rom[574][57] = -8'd9;
        rom[574][58] = -8'd40;
        rom[574][59] = 8'd23;
        rom[574][60] = -8'd31;
        rom[574][61] = -8'd37;
        rom[574][62] = -8'd49;
        rom[574][63] = 8'd3;
        rom[575][0] = 8'd11;
        rom[575][1] = 8'd55;
        rom[575][2] = 8'd22;
        rom[575][3] = -8'd16;
        rom[575][4] = 8'd15;
        rom[575][5] = 8'd19;
        rom[575][6] = 8'd28;
        rom[575][7] = -8'd73;
        rom[575][8] = 8'd24;
        rom[575][9] = 8'd10;
        rom[575][10] = -8'd40;
        rom[575][11] = 8'd15;
        rom[575][12] = -8'd30;
        rom[575][13] = -8'd57;
        rom[575][14] = 8'd31;
        rom[575][15] = 8'd17;
        rom[575][16] = -8'd97;
        rom[575][17] = -8'd15;
        rom[575][18] = -8'd12;
        rom[575][19] = -8'd12;
        rom[575][20] = -8'd11;
        rom[575][21] = 8'd9;
        rom[575][22] = 8'd2;
        rom[575][23] = 8'd3;
        rom[575][24] = -8'd29;
        rom[575][25] = -8'd30;
        rom[575][26] = -8'd21;
        rom[575][27] = 8'd12;
        rom[575][28] = 8'd26;
        rom[575][29] = 8'd37;
        rom[575][30] = 8'd32;
        rom[575][31] = 8'd23;
        rom[575][32] = 8'd27;
        rom[575][33] = 8'd16;
        rom[575][34] = -8'd28;
        rom[575][35] = 8'd11;
        rom[575][36] = 8'd5;
        rom[575][37] = -8'd98;
        rom[575][38] = -8'd8;
        rom[575][39] = 8'd2;
        rom[575][40] = 8'd19;
        rom[575][41] = 8'd35;
        rom[575][42] = 8'd12;
        rom[575][43] = 8'd30;
        rom[575][44] = 8'd16;
        rom[575][45] = -8'd14;
        rom[575][46] = 8'd5;
        rom[575][47] = -8'd30;
        rom[575][48] = -8'd5;
        rom[575][49] = 8'd15;
        rom[575][50] = -8'd20;
        rom[575][51] = 8'd7;
        rom[575][52] = 8'd44;
        rom[575][53] = 8'd37;
        rom[575][54] = 8'd30;
        rom[575][55] = 8'd7;
        rom[575][56] = 8'd8;
        rom[575][57] = -8'd10;
        rom[575][58] = -8'd7;
        rom[575][59] = -8'd22;
        rom[575][60] = 8'd20;
        rom[575][61] = -8'd39;
        rom[575][62] = 8'd16;
        rom[575][63] = 8'd7;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
