module rom_10_dense_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:63][0:9];

    initial begin
        rom[0][0] = -8'd2;
        rom[0][1] = 8'd55;
        rom[0][2] = -8'd6;
        rom[0][3] = -8'd6;
        rom[0][4] = -8'd55;
        rom[0][5] = 8'd30;
        rom[0][6] = -8'd56;
        rom[0][7] = -8'd55;
        rom[0][8] = 8'd58;
        rom[0][9] = 8'd22;
        rom[1][0] = -8'd46;
        rom[1][1] = 8'd4;
        rom[1][2] = 8'd29;
        rom[1][3] = -8'd42;
        rom[1][4] = 8'd36;
        rom[1][5] = -8'd44;
        rom[1][6] = -8'd1;
        rom[1][7] = -8'd41;
        rom[1][8] = 8'd19;
        rom[1][9] = 8'd76;
        rom[2][0] = 8'd0;
        rom[2][1] = 8'd26;
        rom[2][2] = -8'd15;
        rom[2][3] = -8'd36;
        rom[2][4] = 8'd69;
        rom[2][5] = 8'd59;
        rom[2][6] = -8'd1;
        rom[2][7] = 8'd34;
        rom[2][8] = 8'd3;
        rom[2][9] = 8'd9;
        rom[3][0] = 8'd25;
        rom[3][1] = -8'd16;
        rom[3][2] = -8'd28;
        rom[3][3] = 8'd43;
        rom[3][4] = -8'd13;
        rom[3][5] = -8'd45;
        rom[3][6] = -8'd7;
        rom[3][7] = 8'd46;
        rom[3][8] = 8'd57;
        rom[3][9] = 8'd21;
        rom[4][0] = -8'd28;
        rom[4][1] = -8'd19;
        rom[4][2] = -8'd34;
        rom[4][3] = 8'd33;
        rom[4][4] = -8'd32;
        rom[4][5] = 8'd33;
        rom[4][6] = -8'd15;
        rom[4][7] = 8'd69;
        rom[4][8] = -8'd56;
        rom[4][9] = 8'd21;
        rom[5][0] = 8'd13;
        rom[5][1] = -8'd34;
        rom[5][2] = -8'd13;
        rom[5][3] = 8'd42;
        rom[5][4] = -8'd31;
        rom[5][5] = 8'd50;
        rom[5][6] = 8'd37;
        rom[5][7] = 8'd19;
        rom[5][8] = -8'd44;
        rom[5][9] = 8'd1;
        rom[6][0] = -8'd30;
        rom[6][1] = -8'd20;
        rom[6][2] = -8'd24;
        rom[6][3] = -8'd14;
        rom[6][4] = -8'd21;
        rom[6][5] = -8'd7;
        rom[6][6] = 8'd99;
        rom[6][7] = -8'd1;
        rom[6][8] = -8'd10;
        rom[6][9] = -8'd42;
        rom[7][0] = -8'd20;
        rom[7][1] = 8'd15;
        rom[7][2] = -8'd48;
        rom[7][3] = 8'd4;
        rom[7][4] = -8'd20;
        rom[7][5] = 8'd2;
        rom[7][6] = -8'd14;
        rom[7][7] = -8'd10;
        rom[7][8] = 8'd56;
        rom[7][9] = 8'd13;
        rom[8][0] = 8'd33;
        rom[8][1] = -8'd21;
        rom[8][2] = -8'd10;
        rom[8][3] = -8'd17;
        rom[8][4] = 8'd13;
        rom[8][5] = -8'd23;
        rom[8][6] = -8'd46;
        rom[8][7] = 8'd45;
        rom[8][8] = 8'd37;
        rom[8][9] = 8'd15;
        rom[9][0] = 8'd34;
        rom[9][1] = -8'd23;
        rom[9][2] = 8'd15;
        rom[9][3] = -8'd50;
        rom[9][4] = 8'd17;
        rom[9][5] = -8'd42;
        rom[9][6] = -8'd9;
        rom[9][7] = -8'd7;
        rom[9][8] = 8'd24;
        rom[9][9] = -8'd25;
        rom[10][0] = 8'd53;
        rom[10][1] = -8'd43;
        rom[10][2] = 8'd37;
        rom[10][3] = -8'd2;
        rom[10][4] = 8'd14;
        rom[10][5] = 8'd38;
        rom[10][6] = -8'd43;
        rom[10][7] = 8'd14;
        rom[10][8] = -8'd64;
        rom[10][9] = -8'd7;
        rom[11][0] = -8'd57;
        rom[11][1] = -8'd27;
        rom[11][2] = 8'd21;
        rom[11][3] = 8'd40;
        rom[11][4] = -8'd4;
        rom[11][5] = -8'd9;
        rom[11][6] = -8'd15;
        rom[11][7] = 8'd21;
        rom[11][8] = -8'd21;
        rom[11][9] = -8'd53;
        rom[12][0] = 8'd16;
        rom[12][1] = -8'd72;
        rom[12][2] = -8'd6;
        rom[12][3] = -8'd15;
        rom[12][4] = -8'd20;
        rom[12][5] = 8'd31;
        rom[12][6] = 8'd18;
        rom[12][7] = 8'd85;
        rom[12][8] = 8'd46;
        rom[12][9] = -8'd62;
        rom[13][0] = -8'd6;
        rom[13][1] = 8'd3;
        rom[13][2] = -8'd67;
        rom[13][3] = 8'd8;
        rom[13][4] = -8'd12;
        rom[13][5] = 8'd17;
        rom[13][6] = -8'd32;
        rom[13][7] = -8'd15;
        rom[13][8] = -8'd75;
        rom[13][9] = 8'd41;
        rom[14][0] = -8'd25;
        rom[14][1] = -8'd6;
        rom[14][2] = 8'd18;
        rom[14][3] = 8'd9;
        rom[14][4] = -8'd39;
        rom[14][5] = 8'd22;
        rom[14][6] = -8'd62;
        rom[14][7] = -8'd37;
        rom[14][8] = 8'd20;
        rom[14][9] = 8'd44;
        rom[15][0] = 8'd6;
        rom[15][1] = 8'd40;
        rom[15][2] = 8'd3;
        rom[15][3] = -8'd32;
        rom[15][4] = -8'd21;
        rom[15][5] = -8'd36;
        rom[15][6] = -8'd9;
        rom[15][7] = -8'd17;
        rom[15][8] = 8'd58;
        rom[15][9] = 8'd47;
        rom[16][0] = 8'd10;
        rom[16][1] = 8'd19;
        rom[16][2] = -8'd27;
        rom[16][3] = -8'd25;
        rom[16][4] = 8'd22;
        rom[16][5] = -8'd12;
        rom[16][6] = -8'd48;
        rom[16][7] = 8'd66;
        rom[16][8] = -8'd43;
        rom[16][9] = -8'd17;
        rom[17][0] = 8'd20;
        rom[17][1] = -8'd23;
        rom[17][2] = -8'd50;
        rom[17][3] = 8'd9;
        rom[17][4] = -8'd55;
        rom[17][5] = -8'd9;
        rom[17][6] = -8'd4;
        rom[17][7] = -8'd4;
        rom[17][8] = -8'd36;
        rom[17][9] = 8'd14;
        rom[18][0] = -8'd24;
        rom[18][1] = -8'd23;
        rom[18][2] = -8'd42;
        rom[18][3] = 8'd41;
        rom[18][4] = -8'd11;
        rom[18][5] = 8'd26;
        rom[18][6] = -8'd36;
        rom[18][7] = -8'd61;
        rom[18][8] = 8'd22;
        rom[18][9] = -8'd66;
        rom[19][0] = 8'd38;
        rom[19][1] = 8'd43;
        rom[19][2] = -8'd14;
        rom[19][3] = -8'd49;
        rom[19][4] = -8'd66;
        rom[19][5] = -8'd45;
        rom[19][6] = 8'd41;
        rom[19][7] = -8'd10;
        rom[19][8] = -8'd6;
        rom[19][9] = 8'd25;
        rom[20][0] = -8'd17;
        rom[20][1] = -8'd11;
        rom[20][2] = -8'd16;
        rom[20][3] = -8'd27;
        rom[20][4] = 8'd4;
        rom[20][5] = -8'd8;
        rom[20][6] = 8'd21;
        rom[20][7] = -8'd24;
        rom[20][8] = -8'd22;
        rom[20][9] = 8'd25;
        rom[21][0] = -8'd14;
        rom[21][1] = -8'd41;
        rom[21][2] = -8'd11;
        rom[21][3] = -8'd10;
        rom[21][4] = -8'd31;
        rom[21][5] = 8'd24;
        rom[21][6] = 8'd52;
        rom[21][7] = -8'd45;
        rom[21][8] = -8'd26;
        rom[21][9] = -8'd51;
        rom[22][0] = -8'd23;
        rom[22][1] = -8'd25;
        rom[22][2] = 8'd91;
        rom[22][3] = 8'd1;
        rom[22][4] = -8'd18;
        rom[22][5] = 8'd12;
        rom[22][6] = -8'd1;
        rom[22][7] = 8'd41;
        rom[22][8] = -8'd28;
        rom[22][9] = 8'd4;
        rom[23][0] = -8'd28;
        rom[23][1] = 8'd25;
        rom[23][2] = -8'd70;
        rom[23][3] = 8'd5;
        rom[23][4] = 8'd19;
        rom[23][5] = 8'd54;
        rom[23][6] = -8'd28;
        rom[23][7] = 8'd22;
        rom[23][8] = -8'd28;
        rom[23][9] = 8'd44;
        rom[24][0] = -8'd56;
        rom[24][1] = 8'd38;
        rom[24][2] = 8'd45;
        rom[24][3] = 8'd18;
        rom[24][4] = 8'd30;
        rom[24][5] = 8'd41;
        rom[24][6] = -8'd19;
        rom[24][7] = 8'd24;
        rom[24][8] = -8'd54;
        rom[24][9] = -8'd28;
        rom[25][0] = 8'd22;
        rom[25][1] = -8'd26;
        rom[25][2] = -8'd52;
        rom[25][3] = 8'd42;
        rom[25][4] = -8'd66;
        rom[25][5] = -8'd5;
        rom[25][6] = -8'd41;
        rom[25][7] = -8'd7;
        rom[25][8] = 8'd30;
        rom[25][9] = -8'd33;
        rom[26][0] = 8'd38;
        rom[26][1] = -8'd29;
        rom[26][2] = 8'd51;
        rom[26][3] = 8'd5;
        rom[26][4] = -8'd24;
        rom[26][5] = 8'd11;
        rom[26][6] = -8'd47;
        rom[26][7] = -8'd1;
        rom[26][8] = -8'd25;
        rom[26][9] = 8'd20;
        rom[27][0] = 8'd46;
        rom[27][1] = -8'd41;
        rom[27][2] = 8'd2;
        rom[27][3] = 8'd27;
        rom[27][4] = 8'd89;
        rom[27][5] = -8'd3;
        rom[27][6] = -8'd15;
        rom[27][7] = 8'd7;
        rom[27][8] = -8'd88;
        rom[27][9] = -8'd60;
        rom[28][0] = 8'd41;
        rom[28][1] = 8'd15;
        rom[28][2] = 8'd60;
        rom[28][3] = 8'd19;
        rom[28][4] = -8'd17;
        rom[28][5] = -8'd18;
        rom[28][6] = 8'd3;
        rom[28][7] = -8'd13;
        rom[28][8] = 8'd13;
        rom[28][9] = 8'd2;
        rom[29][0] = 8'd21;
        rom[29][1] = 8'd38;
        rom[29][2] = 8'd20;
        rom[29][3] = -8'd8;
        rom[29][4] = -8'd4;
        rom[29][5] = 8'd35;
        rom[29][6] = -8'd66;
        rom[29][7] = -8'd25;
        rom[29][8] = -8'd23;
        rom[29][9] = -8'd32;
        rom[30][0] = -8'd40;
        rom[30][1] = 8'd14;
        rom[30][2] = 8'd49;
        rom[30][3] = 8'd10;
        rom[30][4] = 8'd43;
        rom[30][5] = 8'd19;
        rom[30][6] = -8'd27;
        rom[30][7] = -8'd21;
        rom[30][8] = -8'd75;
        rom[30][9] = -8'd49;
        rom[31][0] = 8'd51;
        rom[31][1] = 8'd14;
        rom[31][2] = -8'd50;
        rom[31][3] = -8'd2;
        rom[31][4] = 8'd45;
        rom[31][5] = 8'd10;
        rom[31][6] = -8'd20;
        rom[31][7] = -8'd31;
        rom[31][8] = 8'd28;
        rom[31][9] = 8'd8;
        rom[32][0] = 8'd17;
        rom[32][1] = 8'd78;
        rom[32][2] = -8'd8;
        rom[32][3] = -8'd34;
        rom[32][4] = -8'd29;
        rom[32][5] = -8'd29;
        rom[32][6] = -8'd13;
        rom[32][7] = 8'd38;
        rom[32][8] = 8'd15;
        rom[32][9] = -8'd7;
        rom[33][0] = -8'd57;
        rom[33][1] = 8'd89;
        rom[33][2] = -8'd31;
        rom[33][3] = 8'd7;
        rom[33][4] = -8'd27;
        rom[33][5] = -8'd8;
        rom[33][6] = -8'd26;
        rom[33][7] = -8'd39;
        rom[33][8] = -8'd60;
        rom[33][9] = 8'd17;
        rom[34][0] = -8'd19;
        rom[34][1] = 8'd46;
        rom[34][2] = -8'd22;
        rom[34][3] = 8'd14;
        rom[34][4] = -8'd40;
        rom[34][5] = 8'd29;
        rom[34][6] = 8'd36;
        rom[34][7] = -8'd16;
        rom[34][8] = 8'd6;
        rom[34][9] = -8'd44;
        rom[35][0] = 8'd35;
        rom[35][1] = -8'd37;
        rom[35][2] = 8'd25;
        rom[35][3] = -8'd10;
        rom[35][4] = -8'd22;
        rom[35][5] = -8'd10;
        rom[35][6] = -8'd51;
        rom[35][7] = 8'd49;
        rom[35][8] = -8'd22;
        rom[35][9] = 8'd13;
        rom[36][0] = -8'd12;
        rom[36][1] = -8'd7;
        rom[36][2] = -8'd8;
        rom[36][3] = 8'd30;
        rom[36][4] = 8'd53;
        rom[36][5] = 8'd5;
        rom[36][6] = -8'd58;
        rom[36][7] = 8'd7;
        rom[36][8] = 8'd32;
        rom[36][9] = -8'd11;
        rom[37][0] = 8'd20;
        rom[37][1] = -8'd20;
        rom[37][2] = 8'd56;
        rom[37][3] = 8'd8;
        rom[37][4] = 8'd32;
        rom[37][5] = -8'd22;
        rom[37][6] = -8'd14;
        rom[37][7] = 8'd13;
        rom[37][8] = -8'd78;
        rom[37][9] = 8'd5;
        rom[38][0] = 8'd10;
        rom[38][1] = -8'd55;
        rom[38][2] = 8'd82;
        rom[38][3] = -8'd18;
        rom[38][4] = -8'd42;
        rom[38][5] = 8'd1;
        rom[38][6] = 8'd7;
        rom[38][7] = -8'd20;
        rom[38][8] = -8'd37;
        rom[38][9] = -8'd51;
        rom[39][0] = -8'd54;
        rom[39][1] = -8'd43;
        rom[39][2] = 8'd27;
        rom[39][3] = 8'd34;
        rom[39][4] = 8'd25;
        rom[39][5] = -8'd2;
        rom[39][6] = 8'd25;
        rom[39][7] = -8'd34;
        rom[39][8] = -8'd37;
        rom[39][9] = -8'd22;
        rom[40][0] = 8'd20;
        rom[40][1] = -8'd7;
        rom[40][2] = -8'd3;
        rom[40][3] = 8'd20;
        rom[40][4] = 8'd36;
        rom[40][5] = 8'd30;
        rom[40][6] = 8'd33;
        rom[40][7] = 8'd27;
        rom[40][8] = -8'd64;
        rom[40][9] = -8'd44;
        rom[41][0] = -8'd34;
        rom[41][1] = -8'd54;
        rom[41][2] = -8'd10;
        rom[41][3] = -8'd20;
        rom[41][4] = 8'd41;
        rom[41][5] = -8'd3;
        rom[41][6] = 8'd37;
        rom[41][7] = 8'd43;
        rom[41][8] = -8'd53;
        rom[41][9] = -8'd53;
        rom[42][0] = -8'd48;
        rom[42][1] = 8'd34;
        rom[42][2] = 8'd15;
        rom[42][3] = 8'd10;
        rom[42][4] = -8'd24;
        rom[42][5] = -8'd34;
        rom[42][6] = 8'd67;
        rom[42][7] = 8'd21;
        rom[42][8] = -8'd10;
        rom[42][9] = 8'd27;
        rom[43][0] = -8'd11;
        rom[43][1] = -8'd19;
        rom[43][2] = 8'd0;
        rom[43][3] = 8'd43;
        rom[43][4] = -8'd24;
        rom[43][5] = 8'd42;
        rom[43][6] = -8'd13;
        rom[43][7] = -8'd22;
        rom[43][8] = -8'd5;
        rom[43][9] = 8'd38;
        rom[44][0] = 8'd34;
        rom[44][1] = -8'd3;
        rom[44][2] = -8'd35;
        rom[44][3] = -8'd18;
        rom[44][4] = -8'd36;
        rom[44][5] = -8'd34;
        rom[44][6] = -8'd55;
        rom[44][7] = 8'd18;
        rom[44][8] = 8'd30;
        rom[44][9] = -8'd12;
        rom[45][0] = -8'd62;
        rom[45][1] = 8'd67;
        rom[45][2] = 8'd12;
        rom[45][3] = 8'd0;
        rom[45][4] = -8'd23;
        rom[45][5] = -8'd6;
        rom[45][6] = 8'd26;
        rom[45][7] = -8'd42;
        rom[45][8] = 8'd42;
        rom[45][9] = 8'd12;
        rom[46][0] = -8'd19;
        rom[46][1] = 8'd42;
        rom[46][2] = -8'd8;
        rom[46][3] = 8'd9;
        rom[46][4] = -8'd6;
        rom[46][5] = -8'd2;
        rom[46][6] = 8'd45;
        rom[46][7] = -8'd43;
        rom[46][8] = -8'd40;
        rom[46][9] = 8'd54;
        rom[47][0] = 8'd27;
        rom[47][1] = 8'd35;
        rom[47][2] = -8'd16;
        rom[47][3] = -8'd3;
        rom[47][4] = -8'd17;
        rom[47][5] = -8'd34;
        rom[47][6] = -8'd1;
        rom[47][7] = -8'd4;
        rom[47][8] = -8'd27;
        rom[47][9] = 8'd69;
        rom[48][0] = -8'd15;
        rom[48][1] = -8'd36;
        rom[48][2] = -8'd5;
        rom[48][3] = -8'd49;
        rom[48][4] = -8'd38;
        rom[48][5] = 8'd92;
        rom[48][6] = -8'd45;
        rom[48][7] = -8'd68;
        rom[48][8] = -8'd15;
        rom[48][9] = -8'd37;
        rom[49][0] = 8'd38;
        rom[49][1] = -8'd56;
        rom[49][2] = 8'd24;
        rom[49][3] = 8'd24;
        rom[49][4] = 8'd34;
        rom[49][5] = 8'd37;
        rom[49][6] = 8'd7;
        rom[49][7] = -8'd35;
        rom[49][8] = 8'd59;
        rom[49][9] = -8'd16;
        rom[50][0] = 8'd4;
        rom[50][1] = 8'd37;
        rom[50][2] = -8'd13;
        rom[50][3] = -8'd3;
        rom[50][4] = 8'd56;
        rom[50][5] = -8'd54;
        rom[50][6] = -8'd40;
        rom[50][7] = -8'd70;
        rom[50][8] = 8'd0;
        rom[50][9] = -8'd5;
        rom[51][0] = -8'd9;
        rom[51][1] = -8'd26;
        rom[51][2] = 8'd6;
        rom[51][3] = -8'd4;
        rom[51][4] = -8'd53;
        rom[51][5] = 8'd44;
        rom[51][6] = 8'd33;
        rom[51][7] = 8'd35;
        rom[51][8] = 8'd28;
        rom[51][9] = -8'd33;
        rom[52][0] = -8'd13;
        rom[52][1] = -8'd98;
        rom[52][2] = 8'd15;
        rom[52][3] = -8'd6;
        rom[52][4] = 8'd36;
        rom[52][5] = -8'd17;
        rom[52][6] = 8'd3;
        rom[52][7] = -8'd8;
        rom[52][8] = 8'd7;
        rom[52][9] = 8'd5;
        rom[53][0] = -8'd30;
        rom[53][1] = -8'd25;
        rom[53][2] = -8'd35;
        rom[53][3] = 8'd61;
        rom[53][4] = 8'd31;
        rom[53][5] = 8'd40;
        rom[53][6] = 8'd17;
        rom[53][7] = 8'd40;
        rom[53][8] = -8'd1;
        rom[53][9] = 8'd7;
        rom[54][0] = -8'd68;
        rom[54][1] = 8'd17;
        rom[54][2] = 8'd42;
        rom[54][3] = -8'd23;
        rom[54][4] = -8'd12;
        rom[54][5] = -8'd25;
        rom[54][6] = 8'd21;
        rom[54][7] = 8'd18;
        rom[54][8] = 8'd39;
        rom[54][9] = -8'd29;
        rom[55][0] = -8'd22;
        rom[55][1] = 8'd30;
        rom[55][2] = -8'd9;
        rom[55][3] = -8'd26;
        rom[55][4] = -8'd26;
        rom[55][5] = 8'd7;
        rom[55][6] = 8'd12;
        rom[55][7] = 8'd38;
        rom[55][8] = 8'd63;
        rom[55][9] = 8'd2;
        rom[56][0] = -8'd26;
        rom[56][1] = -8'd81;
        rom[56][2] = 8'd0;
        rom[56][3] = -8'd2;
        rom[56][4] = 8'd58;
        rom[56][5] = 8'd20;
        rom[56][6] = -8'd20;
        rom[56][7] = 8'd9;
        rom[56][8] = -8'd56;
        rom[56][9] = -8'd55;
        rom[57][0] = 8'd5;
        rom[57][1] = -8'd8;
        rom[57][2] = 8'd15;
        rom[57][3] = -8'd12;
        rom[57][4] = -8'd31;
        rom[57][5] = -8'd19;
        rom[57][6] = 8'd62;
        rom[57][7] = -8'd53;
        rom[57][8] = 8'd35;
        rom[57][9] = 8'd31;
        rom[58][0] = 8'd39;
        rom[58][1] = 8'd29;
        rom[58][2] = 8'd25;
        rom[58][3] = -8'd22;
        rom[58][4] = 8'd33;
        rom[58][5] = -8'd12;
        rom[58][6] = 8'd31;
        rom[58][7] = -8'd56;
        rom[58][8] = -8'd39;
        rom[58][9] = 8'd28;
        rom[59][0] = -8'd71;
        rom[59][1] = 8'd4;
        rom[59][2] = -8'd2;
        rom[59][3] = -8'd13;
        rom[59][4] = 8'd50;
        rom[59][5] = 8'd36;
        rom[59][6] = 8'd17;
        rom[59][7] = 8'd59;
        rom[59][8] = -8'd22;
        rom[59][9] = 8'd33;
        rom[60][0] = 8'd2;
        rom[60][1] = 8'd50;
        rom[60][2] = -8'd30;
        rom[60][3] = -8'd36;
        rom[60][4] = -8'd12;
        rom[60][5] = -8'd31;
        rom[60][6] = 8'd68;
        rom[60][7] = -8'd34;
        rom[60][8] = 8'd17;
        rom[60][9] = 8'd5;
        rom[61][0] = -8'd43;
        rom[61][1] = -8'd16;
        rom[61][2] = -8'd28;
        rom[61][3] = -8'd37;
        rom[61][4] = 8'd13;
        rom[61][5] = -8'd31;
        rom[61][6] = 8'd4;
        rom[61][7] = -8'd12;
        rom[61][8] = 8'd61;
        rom[61][9] = 8'd39;
        rom[62][0] = 8'd29;
        rom[62][1] = -8'd46;
        rom[62][2] = 8'd51;
        rom[62][3] = 8'd6;
        rom[62][4] = 8'd13;
        rom[62][5] = -8'd5;
        rom[62][6] = 8'd22;
        rom[62][7] = -8'd12;
        rom[62][8] = 8'd4;
        rom[62][9] = -8'd68;
        rom[63][0] = 8'd32;
        rom[63][1] = 8'd8;
        rom[63][2] = 8'd33;
        rom[63][3] = 8'd18;
        rom[63][4] = -8'd19;
        rom[63][5] = -8'd42;
        rom[63][6] = 8'd23;
        rom[63][7] = -8'd51;
        rom[63][8] = 8'd30;
        rom[63][9] = -8'd50;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
