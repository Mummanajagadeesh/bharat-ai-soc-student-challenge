module rom_00_conv2d_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:26][0:15];

    initial begin
        rom[0][0] = -8'd23;
        rom[0][1] = -8'd26;
        rom[0][2] = 8'd22;
        rom[0][3] = 8'd25;
        rom[0][4] = 8'd17;
        rom[0][5] = -8'd26;
        rom[0][6] = 8'd19;
        rom[0][7] = -8'd10;
        rom[0][8] = 8'd26;
        rom[0][9] = -8'd11;
        rom[0][10] = 8'd11;
        rom[0][11] = 8'd13;
        rom[0][12] = -8'd1;
        rom[0][13] = 8'd10;
        rom[0][14] = 8'd37;
        rom[0][15] = -8'd11;
        rom[1][0] = -8'd25;
        rom[1][1] = -8'd22;
        rom[1][2] = -8'd12;
        rom[1][3] = 8'd1;
        rom[1][4] = -8'd19;
        rom[1][5] = -8'd8;
        rom[1][6] = 8'd37;
        rom[1][7] = 8'd33;
        rom[1][8] = 8'd8;
        rom[1][9] = -8'd16;
        rom[1][10] = -8'd13;
        rom[1][11] = 8'd5;
        rom[1][12] = 8'd35;
        rom[1][13] = -8'd25;
        rom[1][14] = -8'd4;
        rom[1][15] = -8'd13;
        rom[2][0] = -8'd21;
        rom[2][1] = 8'd7;
        rom[2][2] = 8'd27;
        rom[2][3] = -8'd6;
        rom[2][4] = 8'd13;
        rom[2][5] = 8'd2;
        rom[2][6] = -8'd44;
        rom[2][7] = 8'd6;
        rom[2][8] = 8'd28;
        rom[2][9] = 8'd26;
        rom[2][10] = 8'd28;
        rom[2][11] = -8'd20;
        rom[2][12] = 8'd24;
        rom[2][13] = 8'd11;
        rom[2][14] = -8'd9;
        rom[2][15] = -8'd12;
        rom[3][0] = 8'd0;
        rom[3][1] = -8'd9;
        rom[3][2] = 8'd43;
        rom[3][3] = 8'd33;
        rom[3][4] = -8'd27;
        rom[3][5] = -8'd7;
        rom[3][6] = -8'd14;
        rom[3][7] = -8'd18;
        rom[3][8] = -8'd23;
        rom[3][9] = -8'd17;
        rom[3][10] = -8'd30;
        rom[3][11] = 8'd38;
        rom[3][12] = -8'd2;
        rom[3][13] = 8'd36;
        rom[3][14] = 8'd43;
        rom[3][15] = -8'd24;
        rom[4][0] = 8'd8;
        rom[4][1] = 8'd3;
        rom[4][2] = 8'd21;
        rom[4][3] = 8'd28;
        rom[4][4] = -8'd34;
        rom[4][5] = -8'd14;
        rom[4][6] = 8'd37;
        rom[4][7] = 8'd31;
        rom[4][8] = -8'd34;
        rom[4][9] = -8'd4;
        rom[4][10] = -8'd9;
        rom[4][11] = -8'd20;
        rom[4][12] = -8'd13;
        rom[4][13] = 8'd9;
        rom[4][14] = -8'd28;
        rom[4][15] = 8'd8;
        rom[5][0] = 8'd3;
        rom[5][1] = 8'd13;
        rom[5][2] = 8'd13;
        rom[5][3] = -8'd10;
        rom[5][4] = -8'd28;
        rom[5][5] = 8'd20;
        rom[5][6] = 8'd13;
        rom[5][7] = -8'd36;
        rom[5][8] = -8'd56;
        rom[5][9] = 8'd1;
        rom[5][10] = -8'd3;
        rom[5][11] = -8'd11;
        rom[5][12] = -8'd18;
        rom[5][13] = 8'd33;
        rom[5][14] = -8'd21;
        rom[5][15] = -8'd45;
        rom[6][0] = -8'd4;
        rom[6][1] = -8'd8;
        rom[6][2] = 8'd14;
        rom[6][3] = 8'd11;
        rom[6][4] = 8'd37;
        rom[6][5] = -8'd7;
        rom[6][6] = 8'd4;
        rom[6][7] = -8'd36;
        rom[6][8] = -8'd24;
        rom[6][9] = -8'd4;
        rom[6][10] = -8'd19;
        rom[6][11] = -8'd11;
        rom[6][12] = -8'd20;
        rom[6][13] = 8'd1;
        rom[6][14] = 8'd20;
        rom[6][15] = -8'd24;
        rom[7][0] = -8'd1;
        rom[7][1] = -8'd9;
        rom[7][2] = -8'd9;
        rom[7][3] = 8'd36;
        rom[7][4] = 8'd9;
        rom[7][5] = 8'd11;
        rom[7][6] = -8'd1;
        rom[7][7] = 8'd16;
        rom[7][8] = -8'd19;
        rom[7][9] = -8'd33;
        rom[7][10] = -8'd11;
        rom[7][11] = 8'd0;
        rom[7][12] = 8'd0;
        rom[7][13] = -8'd20;
        rom[7][14] = -8'd37;
        rom[7][15] = 8'd24;
        rom[8][0] = -8'd15;
        rom[8][1] = -8'd8;
        rom[8][2] = 8'd27;
        rom[8][3] = 8'd17;
        rom[8][4] = 8'd7;
        rom[8][5] = 8'd18;
        rom[8][6] = -8'd29;
        rom[8][7] = 8'd9;
        rom[8][8] = -8'd14;
        rom[8][9] = -8'd8;
        rom[8][10] = -8'd44;
        rom[8][11] = 8'd27;
        rom[8][12] = -8'd11;
        rom[8][13] = -8'd11;
        rom[8][14] = -8'd9;
        rom[8][15] = -8'd44;
        rom[9][0] = 8'd2;
        rom[9][1] = -8'd22;
        rom[9][2] = -8'd15;
        rom[9][3] = 8'd53;
        rom[9][4] = -8'd13;
        rom[9][5] = -8'd26;
        rom[9][6] = -8'd17;
        rom[9][7] = -8'd21;
        rom[9][8] = -8'd15;
        rom[9][9] = 8'd12;
        rom[9][10] = -8'd4;
        rom[9][11] = 8'd40;
        rom[9][12] = 8'd39;
        rom[9][13] = -8'd25;
        rom[9][14] = 8'd33;
        rom[9][15] = -8'd10;
        rom[10][0] = 8'd5;
        rom[10][1] = -8'd3;
        rom[10][2] = 8'd11;
        rom[10][3] = 8'd23;
        rom[10][4] = -8'd27;
        rom[10][5] = -8'd1;
        rom[10][6] = 8'd27;
        rom[10][7] = -8'd12;
        rom[10][8] = -8'd49;
        rom[10][9] = -8'd30;
        rom[10][10] = -8'd4;
        rom[10][11] = -8'd8;
        rom[10][12] = 8'd48;
        rom[10][13] = -8'd14;
        rom[10][14] = -8'd16;
        rom[10][15] = -8'd38;
        rom[11][0] = -8'd1;
        rom[11][1] = -8'd24;
        rom[11][2] = 8'd13;
        rom[11][3] = 8'd25;
        rom[11][4] = -8'd14;
        rom[11][5] = 8'd26;
        rom[11][6] = -8'd36;
        rom[11][7] = -8'd5;
        rom[11][8] = -8'd44;
        rom[11][9] = -8'd2;
        rom[11][10] = 8'd27;
        rom[11][11] = -8'd5;
        rom[11][12] = 8'd47;
        rom[11][13] = -8'd32;
        rom[11][14] = 8'd8;
        rom[11][15] = -8'd42;
        rom[12][0] = -8'd24;
        rom[12][1] = 8'd8;
        rom[12][2] = -8'd4;
        rom[12][3] = -8'd73;
        rom[12][4] = 8'd8;
        rom[12][5] = 8'd6;
        rom[12][6] = -8'd28;
        rom[12][7] = -8'd2;
        rom[12][8] = 8'd88;
        rom[12][9] = -8'd13;
        rom[12][10] = -8'd12;
        rom[12][11] = -8'd8;
        rom[12][12] = 8'd26;
        rom[12][13] = 8'd2;
        rom[12][14] = 8'd35;
        rom[12][15] = -8'd42;
        rom[13][0] = -8'd16;
        rom[13][1] = 8'd20;
        rom[13][2] = -8'd3;
        rom[13][3] = -8'd92;
        rom[13][4] = -8'd53;
        rom[13][5] = 8'd20;
        rom[13][6] = 8'd41;
        rom[13][7] = 8'd30;
        rom[13][8] = 8'd95;
        rom[13][9] = -8'd26;
        rom[13][10] = -8'd11;
        rom[13][11] = -8'd55;
        rom[13][12] = 8'd6;
        rom[13][13] = -8'd26;
        rom[13][14] = -8'd51;
        rom[13][15] = 8'd40;
        rom[14][0] = 8'd0;
        rom[14][1] = -8'd8;
        rom[14][2] = 8'd18;
        rom[14][3] = -8'd67;
        rom[14][4] = -8'd7;
        rom[14][5] = 8'd51;
        rom[14][6] = -8'd4;
        rom[14][7] = -8'd38;
        rom[14][8] = 8'd85;
        rom[14][9] = -8'd32;
        rom[14][10] = -8'd8;
        rom[14][11] = 8'd3;
        rom[14][12] = 8'd1;
        rom[14][13] = 8'd4;
        rom[14][14] = -8'd22;
        rom[14][15] = -8'd47;
        rom[15][0] = -8'd15;
        rom[15][1] = -8'd16;
        rom[15][2] = -8'd18;
        rom[15][3] = -8'd2;
        rom[15][4] = 8'd54;
        rom[15][5] = -8'd2;
        rom[15][6] = -8'd32;
        rom[15][7] = 8'd16;
        rom[15][8] = 8'd11;
        rom[15][9] = 8'd36;
        rom[15][10] = -8'd29;
        rom[15][11] = 8'd10;
        rom[15][12] = -8'd19;
        rom[15][13] = 8'd26;
        rom[15][14] = 8'd37;
        rom[15][15] = -8'd32;
        rom[16][0] = -8'd19;
        rom[16][1] = -8'd41;
        rom[16][2] = -8'd27;
        rom[16][3] = -8'd4;
        rom[16][4] = 8'd6;
        rom[16][5] = -8'd29;
        rom[16][6] = 8'd32;
        rom[16][7] = 8'd38;
        rom[16][8] = 8'd15;
        rom[16][9] = -8'd5;
        rom[16][10] = -8'd7;
        rom[16][11] = -8'd21;
        rom[16][12] = -8'd25;
        rom[16][13] = 8'd28;
        rom[16][14] = 8'd3;
        rom[16][15] = 8'd34;
        rom[17][0] = -8'd18;
        rom[17][1] = -8'd26;
        rom[17][2] = 8'd5;
        rom[17][3] = -8'd8;
        rom[17][4] = 8'd11;
        rom[17][5] = 8'd22;
        rom[17][6] = -8'd8;
        rom[17][7] = 8'd0;
        rom[17][8] = 8'd6;
        rom[17][9] = -8'd13;
        rom[17][10] = -8'd21;
        rom[17][11] = -8'd4;
        rom[17][12] = -8'd43;
        rom[17][13] = 8'd27;
        rom[17][14] = 8'd1;
        rom[17][15] = -8'd10;
        rom[18][0] = 8'd6;
        rom[18][1] = 8'd24;
        rom[18][2] = -8'd10;
        rom[18][3] = -8'd12;
        rom[18][4] = -8'd13;
        rom[18][5] = -8'd24;
        rom[18][6] = -8'd9;
        rom[18][7] = -8'd7;
        rom[18][8] = -8'd1;
        rom[18][9] = -8'd15;
        rom[18][10] = -8'd22;
        rom[18][11] = 8'd20;
        rom[18][12] = -8'd9;
        rom[18][13] = 8'd6;
        rom[18][14] = -8'd19;
        rom[18][15] = -8'd15;
        rom[19][0] = -8'd2;
        rom[19][1] = -8'd7;
        rom[19][2] = 8'd5;
        rom[19][3] = -8'd8;
        rom[19][4] = 8'd23;
        rom[19][5] = -8'd13;
        rom[19][6] = 8'd27;
        rom[19][7] = -8'd6;
        rom[19][8] = -8'd21;
        rom[19][9] = -8'd13;
        rom[19][10] = -8'd4;
        rom[19][11] = -8'd32;
        rom[19][12] = -8'd17;
        rom[19][13] = -8'd30;
        rom[19][14] = 8'd20;
        rom[19][15] = -8'd27;
        rom[20][0] = -8'd3;
        rom[20][1] = 8'd24;
        rom[20][2] = -8'd26;
        rom[20][3] = 8'd46;
        rom[20][4] = 8'd36;
        rom[20][5] = 8'd12;
        rom[20][6] = -8'd6;
        rom[20][7] = -8'd38;
        rom[20][8] = 8'd2;
        rom[20][9] = -8'd22;
        rom[20][10] = 8'd25;
        rom[20][11] = 8'd17;
        rom[20][12] = -8'd1;
        rom[20][13] = -8'd12;
        rom[20][14] = 8'd6;
        rom[20][15] = -8'd19;
        rom[21][0] = 8'd3;
        rom[21][1] = 8'd41;
        rom[21][2] = -8'd21;
        rom[21][3] = -8'd29;
        rom[21][4] = 8'd16;
        rom[21][5] = -8'd18;
        rom[21][6] = -8'd26;
        rom[21][7] = 8'd9;
        rom[21][8] = -8'd23;
        rom[21][9] = 8'd14;
        rom[21][10] = 8'd11;
        rom[21][11] = 8'd9;
        rom[21][12] = 8'd5;
        rom[21][13] = -8'd20;
        rom[21][14] = -8'd39;
        rom[21][15] = 8'd2;
        rom[22][0] = 8'd4;
        rom[22][1] = 8'd46;
        rom[22][2] = -8'd28;
        rom[22][3] = -8'd11;
        rom[22][4] = -8'd14;
        rom[22][5] = 8'd11;
        rom[22][6] = -8'd17;
        rom[22][7] = 8'd22;
        rom[22][8] = 8'd2;
        rom[22][9] = -8'd3;
        rom[22][10] = 8'd2;
        rom[22][11] = -8'd33;
        rom[22][12] = -8'd15;
        rom[22][13] = -8'd27;
        rom[22][14] = -8'd35;
        rom[22][15] = 8'd25;
        rom[23][0] = -8'd2;
        rom[23][1] = 8'd41;
        rom[23][2] = -8'd38;
        rom[23][3] = -8'd18;
        rom[23][4] = 8'd43;
        rom[23][5] = 8'd27;
        rom[23][6] = 8'd18;
        rom[23][7] = -8'd28;
        rom[23][8] = -8'd8;
        rom[23][9] = 8'd11;
        rom[23][10] = 8'd38;
        rom[23][11] = 8'd25;
        rom[23][12] = -8'd31;
        rom[23][13] = 8'd10;
        rom[23][14] = 8'd11;
        rom[23][15] = -8'd53;
        rom[24][0] = -8'd1;
        rom[24][1] = 8'd28;
        rom[24][2] = 8'd7;
        rom[24][3] = -8'd8;
        rom[24][4] = 8'd3;
        rom[24][5] = 8'd2;
        rom[24][6] = -8'd12;
        rom[24][7] = 8'd20;
        rom[24][8] = -8'd36;
        rom[24][9] = 8'd6;
        rom[24][10] = 8'd17;
        rom[24][11] = -8'd33;
        rom[24][12] = -8'd7;
        rom[24][13] = 8'd23;
        rom[24][14] = -8'd12;
        rom[24][15] = -8'd26;
        rom[25][0] = -8'd24;
        rom[25][1] = -8'd7;
        rom[25][2] = -8'd4;
        rom[25][3] = 8'd28;
        rom[25][4] = -8'd9;
        rom[25][5] = -8'd21;
        rom[25][6] = -8'd3;
        rom[25][7] = 8'd2;
        rom[25][8] = 8'd8;
        rom[25][9] = 8'd46;
        rom[25][10] = 8'd0;
        rom[25][11] = -8'd3;
        rom[25][12] = -8'd5;
        rom[25][13] = -8'd6;
        rom[25][14] = 8'd30;
        rom[25][15] = 8'd22;
        rom[26][0] = -8'd26;
        rom[26][1] = 8'd4;
        rom[26][2] = -8'd21;
        rom[26][3] = 8'd35;
        rom[26][4] = -8'd17;
        rom[26][5] = -8'd21;
        rom[26][6] = 8'd35;
        rom[26][7] = 8'd16;
        rom[26][8] = -8'd11;
        rom[26][9] = 8'd43;
        rom[26][10] = 8'd20;
        rom[26][11] = 8'd6;
        rom[26][12] = 8'd11;
        rom[26][13] = 8'd33;
        rom[26][14] = 8'd30;
        rom[26][15] = -8'd41;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
