module rom_03_conv2d_2_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:143][0:31];

    initial begin
        rom[0][0] = -8'd6;
        rom[0][1] = -8'd35;
        rom[0][2] = -8'd17;
        rom[0][3] = -8'd16;
        rom[0][4] = -8'd5;
        rom[0][5] = -8'd10;
        rom[0][6] = -8'd13;
        rom[0][7] = 8'd18;
        rom[0][8] = -8'd20;
        rom[0][9] = 8'd10;
        rom[0][10] = -8'd26;
        rom[0][11] = -8'd19;
        rom[0][12] = 8'd4;
        rom[0][13] = 8'd24;
        rom[0][14] = -8'd56;
        rom[0][15] = -8'd20;
        rom[0][16] = 8'd28;
        rom[0][17] = 8'd2;
        rom[0][18] = 8'd11;
        rom[0][19] = 8'd6;
        rom[0][20] = 8'd16;
        rom[0][21] = -8'd3;
        rom[0][22] = 8'd19;
        rom[0][23] = -8'd14;
        rom[0][24] = 8'd29;
        rom[0][25] = -8'd16;
        rom[0][26] = -8'd1;
        rom[0][27] = -8'd30;
        rom[0][28] = 8'd9;
        rom[0][29] = -8'd1;
        rom[0][30] = 8'd9;
        rom[0][31] = -8'd3;
        rom[1][0] = -8'd18;
        rom[1][1] = 8'd12;
        rom[1][2] = -8'd7;
        rom[1][3] = 8'd15;
        rom[1][4] = -8'd20;
        rom[1][5] = -8'd47;
        rom[1][6] = -8'd9;
        rom[1][7] = 8'd0;
        rom[1][8] = 8'd13;
        rom[1][9] = -8'd13;
        rom[1][10] = 8'd30;
        rom[1][11] = -8'd32;
        rom[1][12] = -8'd32;
        rom[1][13] = -8'd11;
        rom[1][14] = -8'd36;
        rom[1][15] = 8'd40;
        rom[1][16] = 8'd3;
        rom[1][17] = -8'd13;
        rom[1][18] = -8'd23;
        rom[1][19] = -8'd2;
        rom[1][20] = -8'd49;
        rom[1][21] = -8'd11;
        rom[1][22] = 8'd5;
        rom[1][23] = -8'd12;
        rom[1][24] = -8'd2;
        rom[1][25] = -8'd27;
        rom[1][26] = -8'd6;
        rom[1][27] = -8'd36;
        rom[1][28] = -8'd42;
        rom[1][29] = -8'd15;
        rom[1][30] = -8'd32;
        rom[1][31] = 8'd16;
        rom[2][0] = 8'd38;
        rom[2][1] = 8'd12;
        rom[2][2] = 8'd13;
        rom[2][3] = 8'd1;
        rom[2][4] = -8'd13;
        rom[2][5] = 8'd19;
        rom[2][6] = -8'd21;
        rom[2][7] = -8'd19;
        rom[2][8] = 8'd13;
        rom[2][9] = 8'd23;
        rom[2][10] = 8'd0;
        rom[2][11] = 8'd24;
        rom[2][12] = 8'd0;
        rom[2][13] = -8'd15;
        rom[2][14] = -8'd4;
        rom[2][15] = 8'd38;
        rom[2][16] = -8'd13;
        rom[2][17] = 8'd0;
        rom[2][18] = 8'd19;
        rom[2][19] = 8'd8;
        rom[2][20] = -8'd22;
        rom[2][21] = -8'd17;
        rom[2][22] = 8'd26;
        rom[2][23] = 8'd4;
        rom[2][24] = -8'd4;
        rom[2][25] = 8'd1;
        rom[2][26] = 8'd6;
        rom[2][27] = -8'd11;
        rom[2][28] = 8'd7;
        rom[2][29] = 8'd8;
        rom[2][30] = -8'd25;
        rom[2][31] = 8'd6;
        rom[3][0] = -8'd5;
        rom[3][1] = 8'd28;
        rom[3][2] = 8'd7;
        rom[3][3] = -8'd2;
        rom[3][4] = 8'd13;
        rom[3][5] = -8'd25;
        rom[3][6] = 8'd8;
        rom[3][7] = 8'd20;
        rom[3][8] = 8'd2;
        rom[3][9] = -8'd2;
        rom[3][10] = -8'd15;
        rom[3][11] = -8'd26;
        rom[3][12] = -8'd16;
        rom[3][13] = -8'd48;
        rom[3][14] = 8'd29;
        rom[3][15] = 8'd37;
        rom[3][16] = 8'd13;
        rom[3][17] = 8'd12;
        rom[3][18] = 8'd14;
        rom[3][19] = -8'd25;
        rom[3][20] = -8'd3;
        rom[3][21] = -8'd13;
        rom[3][22] = -8'd29;
        rom[3][23] = 8'd12;
        rom[3][24] = 8'd12;
        rom[3][25] = -8'd26;
        rom[3][26] = -8'd21;
        rom[3][27] = 8'd14;
        rom[3][28] = -8'd13;
        rom[3][29] = 8'd3;
        rom[3][30] = -8'd19;
        rom[3][31] = -8'd4;
        rom[4][0] = -8'd6;
        rom[4][1] = 8'd6;
        rom[4][2] = -8'd11;
        rom[4][3] = -8'd11;
        rom[4][4] = 8'd14;
        rom[4][5] = 8'd9;
        rom[4][6] = 8'd9;
        rom[4][7] = -8'd2;
        rom[4][8] = 8'd12;
        rom[4][9] = 8'd3;
        rom[4][10] = 8'd26;
        rom[4][11] = -8'd48;
        rom[4][12] = -8'd7;
        rom[4][13] = 8'd2;
        rom[4][14] = -8'd30;
        rom[4][15] = 8'd22;
        rom[4][16] = 8'd12;
        rom[4][17] = -8'd44;
        rom[4][18] = -8'd4;
        rom[4][19] = 8'd4;
        rom[4][20] = 8'd2;
        rom[4][21] = 8'd2;
        rom[4][22] = -8'd4;
        rom[4][23] = -8'd18;
        rom[4][24] = 8'd4;
        rom[4][25] = 8'd14;
        rom[4][26] = -8'd22;
        rom[4][27] = 8'd18;
        rom[4][28] = 8'd9;
        rom[4][29] = -8'd58;
        rom[4][30] = 8'd4;
        rom[4][31] = -8'd4;
        rom[5][0] = 8'd4;
        rom[5][1] = -8'd5;
        rom[5][2] = 8'd36;
        rom[5][3] = 8'd12;
        rom[5][4] = -8'd9;
        rom[5][5] = 8'd36;
        rom[5][6] = 8'd1;
        rom[5][7] = 8'd13;
        rom[5][8] = 8'd17;
        rom[5][9] = 8'd3;
        rom[5][10] = -8'd62;
        rom[5][11] = 8'd0;
        rom[5][12] = 8'd1;
        rom[5][13] = 8'd5;
        rom[5][14] = -8'd3;
        rom[5][15] = 8'd5;
        rom[5][16] = -8'd6;
        rom[5][17] = 8'd3;
        rom[5][18] = -8'd17;
        rom[5][19] = -8'd43;
        rom[5][20] = 8'd9;
        rom[5][21] = 8'd14;
        rom[5][22] = -8'd16;
        rom[5][23] = 8'd12;
        rom[5][24] = 8'd13;
        rom[5][25] = -8'd19;
        rom[5][26] = 8'd18;
        rom[5][27] = -8'd4;
        rom[5][28] = 8'd20;
        rom[5][29] = 8'd2;
        rom[5][30] = 8'd16;
        rom[5][31] = 8'd22;
        rom[6][0] = -8'd38;
        rom[6][1] = 8'd17;
        rom[6][2] = 8'd11;
        rom[6][3] = 8'd1;
        rom[6][4] = 8'd3;
        rom[6][5] = -8'd11;
        rom[6][6] = -8'd18;
        rom[6][7] = 8'd12;
        rom[6][8] = 8'd3;
        rom[6][9] = -8'd2;
        rom[6][10] = 8'd41;
        rom[6][11] = -8'd47;
        rom[6][12] = 8'd10;
        rom[6][13] = 8'd4;
        rom[6][14] = -8'd3;
        rom[6][15] = -8'd40;
        rom[6][16] = -8'd3;
        rom[6][17] = -8'd2;
        rom[6][18] = 8'd1;
        rom[6][19] = 8'd21;
        rom[6][20] = 8'd41;
        rom[6][21] = -8'd11;
        rom[6][22] = 8'd4;
        rom[6][23] = -8'd12;
        rom[6][24] = -8'd55;
        rom[6][25] = -8'd8;
        rom[6][26] = -8'd22;
        rom[6][27] = -8'd18;
        rom[6][28] = 8'd6;
        rom[6][29] = -8'd14;
        rom[6][30] = -8'd48;
        rom[6][31] = 8'd6;
        rom[7][0] = -8'd9;
        rom[7][1] = -8'd12;
        rom[7][2] = 8'd21;
        rom[7][3] = -8'd11;
        rom[7][4] = -8'd14;
        rom[7][5] = 8'd28;
        rom[7][6] = -8'd9;
        rom[7][7] = -8'd27;
        rom[7][8] = 8'd22;
        rom[7][9] = -8'd61;
        rom[7][10] = 8'd24;
        rom[7][11] = 8'd15;
        rom[7][12] = -8'd17;
        rom[7][13] = -8'd9;
        rom[7][14] = -8'd32;
        rom[7][15] = -8'd1;
        rom[7][16] = 8'd0;
        rom[7][17] = -8'd11;
        rom[7][18] = -8'd3;
        rom[7][19] = -8'd2;
        rom[7][20] = -8'd25;
        rom[7][21] = -8'd7;
        rom[7][22] = -8'd6;
        rom[7][23] = 8'd40;
        rom[7][24] = 8'd19;
        rom[7][25] = -8'd22;
        rom[7][26] = -8'd19;
        rom[7][27] = -8'd1;
        rom[7][28] = 8'd7;
        rom[7][29] = 8'd3;
        rom[7][30] = 8'd4;
        rom[7][31] = 8'd1;
        rom[8][0] = 8'd14;
        rom[8][1] = 8'd3;
        rom[8][2] = -8'd17;
        rom[8][3] = -8'd4;
        rom[8][4] = 8'd10;
        rom[8][5] = 8'd36;
        rom[8][6] = 8'd25;
        rom[8][7] = -8'd3;
        rom[8][8] = 8'd11;
        rom[8][9] = -8'd26;
        rom[8][10] = -8'd7;
        rom[8][11] = -8'd12;
        rom[8][12] = 8'd22;
        rom[8][13] = 8'd15;
        rom[8][14] = 8'd4;
        rom[8][15] = 8'd6;
        rom[8][16] = 8'd46;
        rom[8][17] = -8'd24;
        rom[8][18] = 8'd12;
        rom[8][19] = -8'd54;
        rom[8][20] = 8'd17;
        rom[8][21] = 8'd20;
        rom[8][22] = -8'd17;
        rom[8][23] = 8'd11;
        rom[8][24] = -8'd50;
        rom[8][25] = 8'd11;
        rom[8][26] = 8'd12;
        rom[8][27] = 8'd2;
        rom[8][28] = 8'd20;
        rom[8][29] = -8'd39;
        rom[8][30] = 8'd18;
        rom[8][31] = -8'd7;
        rom[9][0] = -8'd26;
        rom[9][1] = -8'd5;
        rom[9][2] = 8'd15;
        rom[9][3] = 8'd18;
        rom[9][4] = -8'd42;
        rom[9][5] = 8'd25;
        rom[9][6] = -8'd12;
        rom[9][7] = 8'd29;
        rom[9][8] = 8'd10;
        rom[9][9] = 8'd5;
        rom[9][10] = 8'd30;
        rom[9][11] = -8'd13;
        rom[9][12] = 8'd11;
        rom[9][13] = -8'd20;
        rom[9][14] = -8'd4;
        rom[9][15] = -8'd1;
        rom[9][16] = 8'd21;
        rom[9][17] = -8'd32;
        rom[9][18] = -8'd5;
        rom[9][19] = 8'd6;
        rom[9][20] = 8'd7;
        rom[9][21] = -8'd25;
        rom[9][22] = -8'd10;
        rom[9][23] = 8'd0;
        rom[9][24] = 8'd8;
        rom[9][25] = 8'd8;
        rom[9][26] = 8'd2;
        rom[9][27] = -8'd13;
        rom[9][28] = -8'd27;
        rom[9][29] = -8'd14;
        rom[9][30] = 8'd31;
        rom[9][31] = -8'd8;
        rom[10][0] = -8'd31;
        rom[10][1] = 8'd41;
        rom[10][2] = 8'd3;
        rom[10][3] = 8'd36;
        rom[10][4] = -8'd11;
        rom[10][5] = -8'd13;
        rom[10][6] = 8'd0;
        rom[10][7] = 8'd3;
        rom[10][8] = -8'd9;
        rom[10][9] = 8'd20;
        rom[10][10] = 8'd15;
        rom[10][11] = 8'd24;
        rom[10][12] = 8'd19;
        rom[10][13] = -8'd2;
        rom[10][14] = 8'd10;
        rom[10][15] = 8'd14;
        rom[10][16] = -8'd20;
        rom[10][17] = -8'd20;
        rom[10][18] = 8'd27;
        rom[10][19] = 8'd23;
        rom[10][20] = -8'd16;
        rom[10][21] = 8'd3;
        rom[10][22] = 8'd54;
        rom[10][23] = -8'd2;
        rom[10][24] = -8'd17;
        rom[10][25] = 8'd30;
        rom[10][26] = -8'd5;
        rom[10][27] = 8'd27;
        rom[10][28] = -8'd7;
        rom[10][29] = -8'd18;
        rom[10][30] = -8'd14;
        rom[10][31] = 8'd9;
        rom[11][0] = 8'd21;
        rom[11][1] = -8'd12;
        rom[11][2] = 8'd41;
        rom[11][3] = -8'd5;
        rom[11][4] = -8'd2;
        rom[11][5] = -8'd2;
        rom[11][6] = -8'd36;
        rom[11][7] = -8'd8;
        rom[11][8] = -8'd15;
        rom[11][9] = 8'd2;
        rom[11][10] = -8'd24;
        rom[11][11] = 8'd3;
        rom[11][12] = -8'd5;
        rom[11][13] = 8'd8;
        rom[11][14] = 8'd11;
        rom[11][15] = 8'd36;
        rom[11][16] = 8'd19;
        rom[11][17] = 8'd5;
        rom[11][18] = -8'd23;
        rom[11][19] = -8'd13;
        rom[11][20] = -8'd15;
        rom[11][21] = 8'd16;
        rom[11][22] = 8'd9;
        rom[11][23] = -8'd28;
        rom[11][24] = 8'd6;
        rom[11][25] = 8'd30;
        rom[11][26] = 8'd9;
        rom[11][27] = 8'd4;
        rom[11][28] = 8'd23;
        rom[11][29] = -8'd11;
        rom[11][30] = -8'd10;
        rom[11][31] = 8'd16;
        rom[12][0] = -8'd24;
        rom[12][1] = 8'd8;
        rom[12][2] = 8'd27;
        rom[12][3] = 8'd31;
        rom[12][4] = -8'd1;
        rom[12][5] = 8'd6;
        rom[12][6] = -8'd6;
        rom[12][7] = 8'd8;
        rom[12][8] = -8'd28;
        rom[12][9] = 8'd17;
        rom[12][10] = 8'd9;
        rom[12][11] = 8'd11;
        rom[12][12] = 8'd22;
        rom[12][13] = -8'd39;
        rom[12][14] = 8'd27;
        rom[12][15] = -8'd4;
        rom[12][16] = -8'd28;
        rom[12][17] = 8'd2;
        rom[12][18] = -8'd3;
        rom[12][19] = -8'd11;
        rom[12][20] = 8'd24;
        rom[12][21] = -8'd10;
        rom[12][22] = -8'd51;
        rom[12][23] = 8'd17;
        rom[12][24] = 8'd12;
        rom[12][25] = -8'd39;
        rom[12][26] = 8'd18;
        rom[12][27] = 8'd3;
        rom[12][28] = -8'd11;
        rom[12][29] = 8'd26;
        rom[12][30] = -8'd13;
        rom[12][31] = 8'd12;
        rom[13][0] = -8'd7;
        rom[13][1] = 8'd6;
        rom[13][2] = 8'd12;
        rom[13][3] = -8'd37;
        rom[13][4] = 8'd21;
        rom[13][5] = 8'd18;
        rom[13][6] = -8'd1;
        rom[13][7] = -8'd4;
        rom[13][8] = 8'd22;
        rom[13][9] = 8'd4;
        rom[13][10] = -8'd17;
        rom[13][11] = -8'd4;
        rom[13][12] = -8'd5;
        rom[13][13] = -8'd3;
        rom[13][14] = -8'd42;
        rom[13][15] = -8'd9;
        rom[13][16] = -8'd2;
        rom[13][17] = 8'd6;
        rom[13][18] = -8'd17;
        rom[13][19] = 8'd28;
        rom[13][20] = -8'd1;
        rom[13][21] = 8'd1;
        rom[13][22] = 8'd43;
        rom[13][23] = 8'd5;
        rom[13][24] = 8'd4;
        rom[13][25] = -8'd3;
        rom[13][26] = -8'd24;
        rom[13][27] = -8'd33;
        rom[13][28] = 8'd10;
        rom[13][29] = 8'd3;
        rom[13][30] = -8'd15;
        rom[13][31] = -8'd6;
        rom[14][0] = -8'd11;
        rom[14][1] = -8'd26;
        rom[14][2] = 8'd25;
        rom[14][3] = 8'd13;
        rom[14][4] = -8'd3;
        rom[14][5] = -8'd13;
        rom[14][6] = 8'd39;
        rom[14][7] = 8'd5;
        rom[14][8] = 8'd16;
        rom[14][9] = -8'd12;
        rom[14][10] = -8'd9;
        rom[14][11] = -8'd7;
        rom[14][12] = 8'd17;
        rom[14][13] = 8'd27;
        rom[14][14] = 8'd5;
        rom[14][15] = 8'd11;
        rom[14][16] = 8'd0;
        rom[14][17] = 8'd20;
        rom[14][18] = 8'd38;
        rom[14][19] = 8'd5;
        rom[14][20] = -8'd33;
        rom[14][21] = -8'd10;
        rom[14][22] = -8'd18;
        rom[14][23] = 8'd8;
        rom[14][24] = 8'd0;
        rom[14][25] = -8'd9;
        rom[14][26] = -8'd16;
        rom[14][27] = -8'd7;
        rom[14][28] = -8'd16;
        rom[14][29] = -8'd58;
        rom[14][30] = 8'd29;
        rom[14][31] = 8'd18;
        rom[15][0] = -8'd19;
        rom[15][1] = 8'd16;
        rom[15][2] = 8'd37;
        rom[15][3] = -8'd14;
        rom[15][4] = 8'd12;
        rom[15][5] = 8'd3;
        rom[15][6] = 8'd8;
        rom[15][7] = -8'd9;
        rom[15][8] = 8'd0;
        rom[15][9] = 8'd23;
        rom[15][10] = 8'd17;
        rom[15][11] = 8'd8;
        rom[15][12] = 8'd8;
        rom[15][13] = -8'd20;
        rom[15][14] = 8'd3;
        rom[15][15] = 8'd14;
        rom[15][16] = -8'd10;
        rom[15][17] = -8'd10;
        rom[15][18] = 8'd5;
        rom[15][19] = 8'd22;
        rom[15][20] = 8'd19;
        rom[15][21] = 8'd7;
        rom[15][22] = 8'd41;
        rom[15][23] = 8'd49;
        rom[15][24] = -8'd20;
        rom[15][25] = 8'd6;
        rom[15][26] = -8'd6;
        rom[15][27] = 8'd0;
        rom[15][28] = 8'd2;
        rom[15][29] = 8'd14;
        rom[15][30] = -8'd39;
        rom[15][31] = 8'd19;
        rom[16][0] = -8'd14;
        rom[16][1] = -8'd34;
        rom[16][2] = -8'd9;
        rom[16][3] = 8'd0;
        rom[16][4] = 8'd15;
        rom[16][5] = -8'd12;
        rom[16][6] = -8'd27;
        rom[16][7] = -8'd29;
        rom[16][8] = -8'd4;
        rom[16][9] = -8'd6;
        rom[16][10] = 8'd9;
        rom[16][11] = -8'd43;
        rom[16][12] = -8'd1;
        rom[16][13] = 8'd4;
        rom[16][14] = -8'd25;
        rom[16][15] = -8'd2;
        rom[16][16] = 8'd20;
        rom[16][17] = -8'd7;
        rom[16][18] = 8'd23;
        rom[16][19] = -8'd17;
        rom[16][20] = 8'd6;
        rom[16][21] = -8'd15;
        rom[16][22] = 8'd5;
        rom[16][23] = -8'd8;
        rom[16][24] = -8'd23;
        rom[16][25] = -8'd26;
        rom[16][26] = 8'd44;
        rom[16][27] = -8'd52;
        rom[16][28] = 8'd18;
        rom[16][29] = -8'd17;
        rom[16][30] = -8'd6;
        rom[16][31] = -8'd10;
        rom[17][0] = 8'd2;
        rom[17][1] = 8'd18;
        rom[17][2] = -8'd10;
        rom[17][3] = 8'd38;
        rom[17][4] = 8'd7;
        rom[17][5] = 8'd4;
        rom[17][6] = -8'd46;
        rom[17][7] = 8'd13;
        rom[17][8] = -8'd16;
        rom[17][9] = 8'd9;
        rom[17][10] = 8'd29;
        rom[17][11] = -8'd42;
        rom[17][12] = -8'd2;
        rom[17][13] = 8'd2;
        rom[17][14] = -8'd54;
        rom[17][15] = 8'd10;
        rom[17][16] = 8'd21;
        rom[17][17] = -8'd23;
        rom[17][18] = -8'd17;
        rom[17][19] = 8'd23;
        rom[17][20] = 8'd15;
        rom[17][21] = -8'd3;
        rom[17][22] = -8'd39;
        rom[17][23] = 8'd0;
        rom[17][24] = 8'd1;
        rom[17][25] = -8'd9;
        rom[17][26] = -8'd12;
        rom[17][27] = -8'd11;
        rom[17][28] = 8'd13;
        rom[17][29] = -8'd28;
        rom[17][30] = -8'd4;
        rom[17][31] = 8'd12;
        rom[18][0] = 8'd35;
        rom[18][1] = 8'd31;
        rom[18][2] = -8'd3;
        rom[18][3] = 8'd22;
        rom[18][4] = -8'd2;
        rom[18][5] = -8'd37;
        rom[18][6] = -8'd42;
        rom[18][7] = 8'd1;
        rom[18][8] = 8'd8;
        rom[18][9] = 8'd21;
        rom[18][10] = 8'd3;
        rom[18][11] = 8'd32;
        rom[18][12] = -8'd57;
        rom[18][13] = 8'd10;
        rom[18][14] = -8'd12;
        rom[18][15] = 8'd6;
        rom[18][16] = -8'd5;
        rom[18][17] = -8'd45;
        rom[18][18] = 8'd44;
        rom[18][19] = 8'd21;
        rom[18][20] = 8'd4;
        rom[18][21] = 8'd6;
        rom[18][22] = 8'd7;
        rom[18][23] = 8'd37;
        rom[18][24] = 8'd3;
        rom[18][25] = -8'd12;
        rom[18][26] = -8'd14;
        rom[18][27] = 8'd1;
        rom[18][28] = -8'd10;
        rom[18][29] = 8'd28;
        rom[18][30] = -8'd28;
        rom[18][31] = -8'd8;
        rom[19][0] = 8'd15;
        rom[19][1] = -8'd14;
        rom[19][2] = 8'd19;
        rom[19][3] = 8'd34;
        rom[19][4] = 8'd3;
        rom[19][5] = 8'd1;
        rom[19][6] = -8'd20;
        rom[19][7] = 8'd1;
        rom[19][8] = -8'd6;
        rom[19][9] = 8'd22;
        rom[19][10] = -8'd6;
        rom[19][11] = -8'd10;
        rom[19][12] = 8'd3;
        rom[19][13] = -8'd19;
        rom[19][14] = 8'd0;
        rom[19][15] = 8'd57;
        rom[19][16] = 8'd13;
        rom[19][17] = -8'd19;
        rom[19][18] = 8'd31;
        rom[19][19] = -8'd7;
        rom[19][20] = -8'd11;
        rom[19][21] = -8'd2;
        rom[19][22] = -8'd49;
        rom[19][23] = -8'd41;
        rom[19][24] = 8'd19;
        rom[19][25] = 8'd12;
        rom[19][26] = -8'd13;
        rom[19][27] = 8'd8;
        rom[19][28] = 8'd16;
        rom[19][29] = -8'd55;
        rom[19][30] = 8'd26;
        rom[19][31] = -8'd5;
        rom[20][0] = 8'd7;
        rom[20][1] = -8'd9;
        rom[20][2] = 8'd7;
        rom[20][3] = 8'd8;
        rom[20][4] = 8'd14;
        rom[20][5] = 8'd6;
        rom[20][6] = -8'd13;
        rom[20][7] = 8'd11;
        rom[20][8] = 8'd13;
        rom[20][9] = -8'd9;
        rom[20][10] = 8'd12;
        rom[20][11] = -8'd2;
        rom[20][12] = 8'd10;
        rom[20][13] = 8'd39;
        rom[20][14] = -8'd9;
        rom[20][15] = 8'd26;
        rom[20][16] = 8'd18;
        rom[20][17] = -8'd50;
        rom[20][18] = 8'd1;
        rom[20][19] = -8'd16;
        rom[20][20] = -8'd17;
        rom[20][21] = -8'd13;
        rom[20][22] = -8'd16;
        rom[20][23] = -8'd3;
        rom[20][24] = -8'd25;
        rom[20][25] = -8'd9;
        rom[20][26] = 8'd12;
        rom[20][27] = 8'd23;
        rom[20][28] = 8'd18;
        rom[20][29] = -8'd79;
        rom[20][30] = 8'd5;
        rom[20][31] = 8'd15;
        rom[21][0] = 8'd7;
        rom[21][1] = -8'd4;
        rom[21][2] = 8'd22;
        rom[21][3] = -8'd25;
        rom[21][4] = 8'd9;
        rom[21][5] = 8'd21;
        rom[21][6] = 8'd33;
        rom[21][7] = -8'd18;
        rom[21][8] = 8'd11;
        rom[21][9] = -8'd22;
        rom[21][10] = -8'd21;
        rom[21][11] = 8'd20;
        rom[21][12] = -8'd18;
        rom[21][13] = -8'd22;
        rom[21][14] = 8'd7;
        rom[21][15] = 8'd34;
        rom[21][16] = -8'd5;
        rom[21][17] = 8'd3;
        rom[21][18] = -8'd5;
        rom[21][19] = -8'd26;
        rom[21][20] = -8'd14;
        rom[21][21] = 8'd6;
        rom[21][22] = -8'd44;
        rom[21][23] = 8'd13;
        rom[21][24] = 8'd8;
        rom[21][25] = 8'd13;
        rom[21][26] = 8'd25;
        rom[21][27] = -8'd14;
        rom[21][28] = -8'd48;
        rom[21][29] = -8'd2;
        rom[21][30] = -8'd13;
        rom[21][31] = 8'd30;
        rom[22][0] = -8'd40;
        rom[22][1] = -8'd8;
        rom[22][2] = -8'd6;
        rom[22][3] = 8'd46;
        rom[22][4] = -8'd5;
        rom[22][5] = -8'd75;
        rom[22][6] = -8'd58;
        rom[22][7] = -8'd10;
        rom[22][8] = -8'd5;
        rom[22][9] = 8'd8;
        rom[22][10] = -8'd8;
        rom[22][11] = -8'd17;
        rom[22][12] = 8'd3;
        rom[22][13] = 8'd29;
        rom[22][14] = -8'd11;
        rom[22][15] = -8'd44;
        rom[22][16] = 8'd19;
        rom[22][17] = -8'd5;
        rom[22][18] = 8'd7;
        rom[22][19] = 8'd21;
        rom[22][20] = 8'd40;
        rom[22][21] = -8'd16;
        rom[22][22] = 8'd1;
        rom[22][23] = -8'd9;
        rom[22][24] = -8'd61;
        rom[22][25] = -8'd65;
        rom[22][26] = -8'd3;
        rom[22][27] = -8'd11;
        rom[22][28] = 8'd14;
        rom[22][29] = 8'd0;
        rom[22][30] = 8'd15;
        rom[22][31] = 8'd7;
        rom[23][0] = -8'd37;
        rom[23][1] = -8'd17;
        rom[23][2] = 8'd14;
        rom[23][3] = -8'd39;
        rom[23][4] = 8'd9;
        rom[23][5] = 8'd21;
        rom[23][6] = 8'd15;
        rom[23][7] = -8'd17;
        rom[23][8] = 8'd10;
        rom[23][9] = -8'd31;
        rom[23][10] = 8'd36;
        rom[23][11] = 8'd25;
        rom[23][12] = -8'd20;
        rom[23][13] = -8'd29;
        rom[23][14] = -8'd23;
        rom[23][15] = -8'd17;
        rom[23][16] = -8'd7;
        rom[23][17] = 8'd1;
        rom[23][18] = 8'd2;
        rom[23][19] = 8'd8;
        rom[23][20] = 8'd24;
        rom[23][21] = 8'd2;
        rom[23][22] = -8'd19;
        rom[23][23] = 8'd32;
        rom[23][24] = 8'd9;
        rom[23][25] = 8'd24;
        rom[23][26] = 8'd17;
        rom[23][27] = 8'd12;
        rom[23][28] = -8'd18;
        rom[23][29] = -8'd19;
        rom[23][30] = -8'd27;
        rom[23][31] = 8'd19;
        rom[24][0] = -8'd6;
        rom[24][1] = -8'd22;
        rom[24][2] = -8'd1;
        rom[24][3] = -8'd5;
        rom[24][4] = 8'd13;
        rom[24][5] = 8'd3;
        rom[24][6] = 8'd22;
        rom[24][7] = 8'd4;
        rom[24][8] = 8'd36;
        rom[24][9] = -8'd8;
        rom[24][10] = -8'd20;
        rom[24][11] = 8'd27;
        rom[24][12] = -8'd25;
        rom[24][13] = 8'd23;
        rom[24][14] = -8'd1;
        rom[24][15] = -8'd12;
        rom[24][16] = 8'd18;
        rom[24][17] = -8'd4;
        rom[24][18] = 8'd16;
        rom[24][19] = -8'd42;
        rom[24][20] = 8'd30;
        rom[24][21] = 8'd23;
        rom[24][22] = -8'd13;
        rom[24][23] = 8'd21;
        rom[24][24] = -8'd125;
        rom[24][25] = -8'd9;
        rom[24][26] = 8'd19;
        rom[24][27] = -8'd22;
        rom[24][28] = 8'd5;
        rom[24][29] = -8'd28;
        rom[24][30] = -8'd4;
        rom[24][31] = -8'd9;
        rom[25][0] = -8'd18;
        rom[25][1] = -8'd16;
        rom[25][2] = 8'd14;
        rom[25][3] = 8'd29;
        rom[25][4] = -8'd1;
        rom[25][5] = 8'd16;
        rom[25][6] = 8'd9;
        rom[25][7] = 8'd18;
        rom[25][8] = 8'd4;
        rom[25][9] = -8'd2;
        rom[25][10] = 8'd16;
        rom[25][11] = -8'd20;
        rom[25][12] = 8'd35;
        rom[25][13] = -8'd14;
        rom[25][14] = 8'd7;
        rom[25][15] = 8'd28;
        rom[25][16] = 8'd10;
        rom[25][17] = -8'd1;
        rom[25][18] = -8'd28;
        rom[25][19] = -8'd24;
        rom[25][20] = -8'd9;
        rom[25][21] = -8'd40;
        rom[25][22] = -8'd16;
        rom[25][23] = -8'd3;
        rom[25][24] = -8'd45;
        rom[25][25] = -8'd51;
        rom[25][26] = -8'd10;
        rom[25][27] = -8'd37;
        rom[25][28] = -8'd37;
        rom[25][29] = -8'd49;
        rom[25][30] = 8'd37;
        rom[25][31] = 8'd4;
        rom[26][0] = -8'd64;
        rom[26][1] = 8'd40;
        rom[26][2] = 8'd18;
        rom[26][3] = 8'd26;
        rom[26][4] = 8'd16;
        rom[26][5] = -8'd79;
        rom[26][6] = -8'd15;
        rom[26][7] = 8'd15;
        rom[26][8] = -8'd11;
        rom[26][9] = 8'd5;
        rom[26][10] = 8'd3;
        rom[26][11] = 8'd19;
        rom[26][12] = 8'd16;
        rom[26][13] = 8'd11;
        rom[26][14] = -8'd8;
        rom[26][15] = 8'd1;
        rom[26][16] = 8'd13;
        rom[26][17] = -8'd43;
        rom[26][18] = 8'd24;
        rom[26][19] = 8'd44;
        rom[26][20] = -8'd5;
        rom[26][21] = -8'd35;
        rom[26][22] = 8'd8;
        rom[26][23] = 8'd30;
        rom[26][24] = -8'd19;
        rom[26][25] = -8'd11;
        rom[26][26] = 8'd23;
        rom[26][27] = 8'd12;
        rom[26][28] = 8'd21;
        rom[26][29] = -8'd13;
        rom[26][30] = -8'd21;
        rom[26][31] = 8'd5;
        rom[27][0] = 8'd1;
        rom[27][1] = -8'd20;
        rom[27][2] = 8'd7;
        rom[27][3] = -8'd8;
        rom[27][4] = 8'd2;
        rom[27][5] = 8'd1;
        rom[27][6] = -8'd9;
        rom[27][7] = 8'd8;
        rom[27][8] = -8'd7;
        rom[27][9] = 8'd11;
        rom[27][10] = -8'd4;
        rom[27][11] = -8'd9;
        rom[27][12] = -8'd18;
        rom[27][13] = 8'd5;
        rom[27][14] = 8'd11;
        rom[27][15] = 8'd19;
        rom[27][16] = -8'd9;
        rom[27][17] = 8'd7;
        rom[27][18] = -8'd10;
        rom[27][19] = -8'd7;
        rom[27][20] = -8'd22;
        rom[27][21] = 8'd10;
        rom[27][22] = -8'd24;
        rom[27][23] = -8'd4;
        rom[27][24] = 8'd14;
        rom[27][25] = 8'd14;
        rom[27][26] = -8'd11;
        rom[27][27] = -8'd2;
        rom[27][28] = -8'd24;
        rom[27][29] = -8'd41;
        rom[27][30] = 8'd3;
        rom[27][31] = 8'd45;
        rom[28][0] = -8'd2;
        rom[28][1] = -8'd4;
        rom[28][2] = 8'd37;
        rom[28][3] = -8'd18;
        rom[28][4] = 8'd19;
        rom[28][5] = 8'd55;
        rom[28][6] = -8'd14;
        rom[28][7] = 8'd15;
        rom[28][8] = -8'd10;
        rom[28][9] = 8'd40;
        rom[28][10] = 8'd26;
        rom[28][11] = 8'd29;
        rom[28][12] = -8'd2;
        rom[28][13] = -8'd16;
        rom[28][14] = 8'd4;
        rom[28][15] = -8'd1;
        rom[28][16] = 8'd7;
        rom[28][17] = -8'd2;
        rom[28][18] = -8'd25;
        rom[28][19] = -8'd9;
        rom[28][20] = 8'd2;
        rom[28][21] = 8'd8;
        rom[28][22] = -8'd45;
        rom[28][23] = -8'd2;
        rom[28][24] = 8'd10;
        rom[28][25] = -8'd29;
        rom[28][26] = 8'd18;
        rom[28][27] = -8'd8;
        rom[28][28] = -8'd12;
        rom[28][29] = 8'd40;
        rom[28][30] = 8'd21;
        rom[28][31] = -8'd2;
        rom[29][0] = -8'd29;
        rom[29][1] = 8'd9;
        rom[29][2] = 8'd8;
        rom[29][3] = -8'd29;
        rom[29][4] = 8'd39;
        rom[29][5] = -8'd2;
        rom[29][6] = 8'd17;
        rom[29][7] = -8'd5;
        rom[29][8] = -8'd7;
        rom[29][9] = 8'd23;
        rom[29][10] = -8'd36;
        rom[29][11] = -8'd12;
        rom[29][12] = -8'd29;
        rom[29][13] = 8'd4;
        rom[29][14] = -8'd41;
        rom[29][15] = 8'd10;
        rom[29][16] = -8'd7;
        rom[29][17] = 8'd5;
        rom[29][18] = 8'd14;
        rom[29][19] = 8'd4;
        rom[29][20] = -8'd35;
        rom[29][21] = 8'd9;
        rom[29][22] = 8'd15;
        rom[29][23] = 8'd15;
        rom[29][24] = 8'd11;
        rom[29][25] = -8'd28;
        rom[29][26] = -8'd1;
        rom[29][27] = -8'd14;
        rom[29][28] = -8'd44;
        rom[29][29] = 8'd19;
        rom[29][30] = -8'd11;
        rom[29][31] = -8'd17;
        rom[30][0] = -8'd12;
        rom[30][1] = 8'd13;
        rom[30][2] = 8'd11;
        rom[30][3] = 8'd30;
        rom[30][4] = 8'd14;
        rom[30][5] = 8'd14;
        rom[30][6] = 8'd36;
        rom[30][7] = -8'd5;
        rom[30][8] = -8'd25;
        rom[30][9] = 8'd14;
        rom[30][10] = -8'd22;
        rom[30][11] = -8'd23;
        rom[30][12] = 8'd19;
        rom[30][13] = 8'd13;
        rom[30][14] = -8'd42;
        rom[30][15] = -8'd1;
        rom[30][16] = 8'd23;
        rom[30][17] = -8'd2;
        rom[30][18] = 8'd24;
        rom[30][19] = -8'd7;
        rom[30][20] = -8'd28;
        rom[30][21] = 8'd35;
        rom[30][22] = -8'd27;
        rom[30][23] = 8'd7;
        rom[30][24] = 8'd18;
        rom[30][25] = -8'd8;
        rom[30][26] = 8'd1;
        rom[30][27] = 8'd9;
        rom[30][28] = -8'd14;
        rom[30][29] = -8'd61;
        rom[30][30] = 8'd6;
        rom[30][31] = 8'd24;
        rom[31][0] = -8'd49;
        rom[31][1] = 8'd18;
        rom[31][2] = 8'd6;
        rom[31][3] = -8'd13;
        rom[31][4] = 8'd24;
        rom[31][5] = -8'd50;
        rom[31][6] = 8'd7;
        rom[31][7] = 8'd23;
        rom[31][8] = -8'd11;
        rom[31][9] = -8'd32;
        rom[31][10] = 8'd18;
        rom[31][11] = -8'd11;
        rom[31][12] = 8'd1;
        rom[31][13] = -8'd50;
        rom[31][14] = -8'd7;
        rom[31][15] = -8'd18;
        rom[31][16] = 8'd17;
        rom[31][17] = -8'd2;
        rom[31][18] = -8'd2;
        rom[31][19] = 8'd30;
        rom[31][20] = 8'd0;
        rom[31][21] = 8'd15;
        rom[31][22] = -8'd5;
        rom[31][23] = 8'd38;
        rom[31][24] = 8'd0;
        rom[31][25] = -8'd21;
        rom[31][26] = -8'd13;
        rom[31][27] = 8'd5;
        rom[31][28] = -8'd23;
        rom[31][29] = 8'd1;
        rom[31][30] = -8'd25;
        rom[31][31] = 8'd30;
        rom[32][0] = -8'd53;
        rom[32][1] = -8'd6;
        rom[32][2] = 8'd5;
        rom[32][3] = -8'd6;
        rom[32][4] = -8'd26;
        rom[32][5] = -8'd26;
        rom[32][6] = -8'd63;
        rom[32][7] = -8'd11;
        rom[32][8] = 8'd11;
        rom[32][9] = -8'd8;
        rom[32][10] = 8'd22;
        rom[32][11] = 8'd7;
        rom[32][12] = -8'd17;
        rom[32][13] = 8'd7;
        rom[32][14] = -8'd30;
        rom[32][15] = -8'd47;
        rom[32][16] = 8'd8;
        rom[32][17] = 8'd26;
        rom[32][18] = -8'd22;
        rom[32][19] = 8'd15;
        rom[32][20] = 8'd45;
        rom[32][21] = 8'd30;
        rom[32][22] = 8'd8;
        rom[32][23] = -8'd1;
        rom[32][24] = -8'd5;
        rom[32][25] = -8'd27;
        rom[32][26] = -8'd7;
        rom[32][27] = -8'd5;
        rom[32][28] = -8'd9;
        rom[32][29] = 8'd31;
        rom[32][30] = -8'd29;
        rom[32][31] = -8'd18;
        rom[33][0] = -8'd1;
        rom[33][1] = 8'd22;
        rom[33][2] = -8'd18;
        rom[33][3] = 8'd20;
        rom[33][4] = -8'd21;
        rom[33][5] = 8'd4;
        rom[33][6] = -8'd34;
        rom[33][7] = 8'd11;
        rom[33][8] = -8'd4;
        rom[33][9] = -8'd25;
        rom[33][10] = 8'd19;
        rom[33][11] = -8'd1;
        rom[33][12] = 8'd15;
        rom[33][13] = -8'd27;
        rom[33][14] = -8'd13;
        rom[33][15] = -8'd31;
        rom[33][16] = -8'd12;
        rom[33][17] = -8'd30;
        rom[33][18] = -8'd11;
        rom[33][19] = -8'd4;
        rom[33][20] = 8'd18;
        rom[33][21] = 8'd11;
        rom[33][22] = -8'd40;
        rom[33][23] = 8'd7;
        rom[33][24] = 8'd11;
        rom[33][25] = -8'd49;
        rom[33][26] = 8'd15;
        rom[33][27] = 8'd25;
        rom[33][28] = 8'd15;
        rom[33][29] = -8'd46;
        rom[33][30] = 8'd25;
        rom[33][31] = 8'd14;
        rom[34][0] = 8'd28;
        rom[34][1] = -8'd15;
        rom[34][2] = 8'd23;
        rom[34][3] = 8'd2;
        rom[34][4] = -8'd1;
        rom[34][5] = -8'd24;
        rom[34][6] = -8'd48;
        rom[34][7] = 8'd7;
        rom[34][8] = -8'd7;
        rom[34][9] = 8'd3;
        rom[34][10] = -8'd1;
        rom[34][11] = 8'd16;
        rom[34][12] = -8'd45;
        rom[34][13] = 8'd17;
        rom[34][14] = -8'd1;
        rom[34][15] = -8'd26;
        rom[34][16] = -8'd8;
        rom[34][17] = -8'd53;
        rom[34][18] = 8'd4;
        rom[34][19] = -8'd12;
        rom[34][20] = 8'd26;
        rom[34][21] = -8'd29;
        rom[34][22] = -8'd33;
        rom[34][23] = 8'd12;
        rom[34][24] = 8'd12;
        rom[34][25] = 8'd11;
        rom[34][26] = 8'd47;
        rom[34][27] = -8'd16;
        rom[34][28] = 8'd47;
        rom[34][29] = 8'd22;
        rom[34][30] = 8'd19;
        rom[34][31] = -8'd14;
        rom[35][0] = -8'd1;
        rom[35][1] = -8'd54;
        rom[35][2] = 8'd0;
        rom[35][3] = 8'd28;
        rom[35][4] = -8'd32;
        rom[35][5] = -8'd18;
        rom[35][6] = -8'd1;
        rom[35][7] = 8'd9;
        rom[35][8] = -8'd39;
        rom[35][9] = -8'd10;
        rom[35][10] = 8'd13;
        rom[35][11] = 8'd10;
        rom[35][12] = 8'd28;
        rom[35][13] = -8'd57;
        rom[35][14] = -8'd18;
        rom[35][15] = 8'd38;
        rom[35][16] = 8'd23;
        rom[35][17] = 8'd4;
        rom[35][18] = 8'd1;
        rom[35][19] = -8'd3;
        rom[35][20] = 8'd0;
        rom[35][21] = 8'd6;
        rom[35][22] = -8'd13;
        rom[35][23] = -8'd33;
        rom[35][24] = -8'd12;
        rom[35][25] = -8'd4;
        rom[35][26] = -8'd26;
        rom[35][27] = -8'd3;
        rom[35][28] = 8'd16;
        rom[35][29] = -8'd34;
        rom[35][30] = 8'd14;
        rom[35][31] = 8'd8;
        rom[36][0] = 8'd14;
        rom[36][1] = -8'd16;
        rom[36][2] = -8'd7;
        rom[36][3] = 8'd9;
        rom[36][4] = -8'd19;
        rom[36][5] = 8'd1;
        rom[36][6] = -8'd4;
        rom[36][7] = -8'd13;
        rom[36][8] = -8'd10;
        rom[36][9] = 8'd4;
        rom[36][10] = -8'd21;
        rom[36][11] = 8'd42;
        rom[36][12] = 8'd6;
        rom[36][13] = 8'd20;
        rom[36][14] = 8'd0;
        rom[36][15] = 8'd2;
        rom[36][16] = 8'd17;
        rom[36][17] = 8'd3;
        rom[36][18] = -8'd15;
        rom[36][19] = 8'd12;
        rom[36][20] = 8'd19;
        rom[36][21] = 8'd23;
        rom[36][22] = -8'd2;
        rom[36][23] = -8'd19;
        rom[36][24] = -8'd9;
        rom[36][25] = -8'd34;
        rom[36][26] = -8'd15;
        rom[36][27] = 8'd20;
        rom[36][28] = 8'd4;
        rom[36][29] = -8'd72;
        rom[36][30] = -8'd10;
        rom[36][31] = -8'd7;
        rom[37][0] = 8'd31;
        rom[37][1] = -8'd23;
        rom[37][2] = -8'd21;
        rom[37][3] = 8'd11;
        rom[37][4] = -8'd17;
        rom[37][5] = 8'd1;
        rom[37][6] = 8'd26;
        rom[37][7] = -8'd12;
        rom[37][8] = 8'd2;
        rom[37][9] = -8'd16;
        rom[37][10] = 8'd26;
        rom[37][11] = 8'd6;
        rom[37][12] = -8'd10;
        rom[37][13] = 8'd15;
        rom[37][14] = 8'd18;
        rom[37][15] = 8'd22;
        rom[37][16] = -8'd34;
        rom[37][17] = 8'd14;
        rom[37][18] = 8'd6;
        rom[37][19] = -8'd1;
        rom[37][20] = 8'd13;
        rom[37][21] = -8'd16;
        rom[37][22] = -8'd7;
        rom[37][23] = 8'd19;
        rom[37][24] = 8'd9;
        rom[37][25] = 8'd33;
        rom[37][26] = 8'd18;
        rom[37][27] = 8'd2;
        rom[37][28] = 8'd12;
        rom[37][29] = -8'd6;
        rom[37][30] = -8'd47;
        rom[37][31] = 8'd47;
        rom[38][0] = -8'd4;
        rom[38][1] = 8'd5;
        rom[38][2] = 8'd17;
        rom[38][3] = 8'd34;
        rom[38][4] = -8'd7;
        rom[38][5] = -8'd86;
        rom[38][6] = -8'd6;
        rom[38][7] = 8'd6;
        rom[38][8] = 8'd5;
        rom[38][9] = 8'd11;
        rom[38][10] = -8'd48;
        rom[38][11] = 8'd6;
        rom[38][12] = 8'd16;
        rom[38][13] = 8'd21;
        rom[38][14] = 8'd9;
        rom[38][15] = -8'd34;
        rom[38][16] = 8'd20;
        rom[38][17] = -8'd18;
        rom[38][18] = 8'd10;
        rom[38][19] = -8'd15;
        rom[38][20] = 8'd40;
        rom[38][21] = 8'd13;
        rom[38][22] = -8'd8;
        rom[38][23] = 8'd14;
        rom[38][24] = 8'd31;
        rom[38][25] = -8'd54;
        rom[38][26] = 8'd18;
        rom[38][27] = 8'd0;
        rom[38][28] = 8'd25;
        rom[38][29] = 8'd14;
        rom[38][30] = 8'd17;
        rom[38][31] = 8'd0;
        rom[39][0] = 8'd4;
        rom[39][1] = -8'd37;
        rom[39][2] = 8'd14;
        rom[39][3] = -8'd25;
        rom[39][4] = 8'd4;
        rom[39][5] = -8'd15;
        rom[39][6] = 8'd11;
        rom[39][7] = -8'd10;
        rom[39][8] = 8'd9;
        rom[39][9] = -8'd6;
        rom[39][10] = 8'd39;
        rom[39][11] = 8'd2;
        rom[39][12] = -8'd36;
        rom[39][13] = -8'd21;
        rom[39][14] = -8'd1;
        rom[39][15] = -8'd16;
        rom[39][16] = -8'd5;
        rom[39][17] = 8'd40;
        rom[39][18] = 8'd17;
        rom[39][19] = 8'd22;
        rom[39][20] = 8'd28;
        rom[39][21] = -8'd28;
        rom[39][22] = 8'd11;
        rom[39][23] = 8'd27;
        rom[39][24] = -8'd17;
        rom[39][25] = 8'd24;
        rom[39][26] = -8'd10;
        rom[39][27] = 8'd4;
        rom[39][28] = -8'd11;
        rom[39][29] = -8'd6;
        rom[39][30] = -8'd28;
        rom[39][31] = 8'd27;
        rom[40][0] = -8'd1;
        rom[40][1] = -8'd11;
        rom[40][2] = 8'd8;
        rom[40][3] = 8'd19;
        rom[40][4] = -8'd3;
        rom[40][5] = -8'd26;
        rom[40][6] = 8'd4;
        rom[40][7] = -8'd15;
        rom[40][8] = 8'd16;
        rom[40][9] = 8'd14;
        rom[40][10] = -8'd3;
        rom[40][11] = 8'd15;
        rom[40][12] = -8'd14;
        rom[40][13] = 8'd35;
        rom[40][14] = -8'd10;
        rom[40][15] = -8'd6;
        rom[40][16] = -8'd15;
        rom[40][17] = 8'd21;
        rom[40][18] = 8'd7;
        rom[40][19] = -8'd3;
        rom[40][20] = 8'd22;
        rom[40][21] = 8'd39;
        rom[40][22] = 8'd17;
        rom[40][23] = 8'd16;
        rom[40][24] = 8'd0;
        rom[40][25] = -8'd33;
        rom[40][26] = -8'd2;
        rom[40][27] = -8'd7;
        rom[40][28] = 8'd10;
        rom[40][29] = -8'd20;
        rom[40][30] = -8'd12;
        rom[40][31] = 8'd9;
        rom[41][0] = -8'd16;
        rom[41][1] = 8'd47;
        rom[41][2] = -8'd12;
        rom[41][3] = 8'd43;
        rom[41][4] = 8'd57;
        rom[41][5] = 8'd17;
        rom[41][6] = 8'd18;
        rom[41][7] = 8'd0;
        rom[41][8] = 8'd33;
        rom[41][9] = 8'd14;
        rom[41][10] = -8'd24;
        rom[41][11] = 8'd28;
        rom[41][12] = 8'd37;
        rom[41][13] = -8'd32;
        rom[41][14] = 8'd16;
        rom[41][15] = 8'd21;
        rom[41][16] = 8'd8;
        rom[41][17] = -8'd2;
        rom[41][18] = -8'd9;
        rom[41][19] = 8'd10;
        rom[41][20] = -8'd27;
        rom[41][21] = -8'd6;
        rom[41][22] = -8'd4;
        rom[41][23] = -8'd17;
        rom[41][24] = 8'd16;
        rom[41][25] = -8'd37;
        rom[41][26] = -8'd21;
        rom[41][27] = -8'd11;
        rom[41][28] = -8'd47;
        rom[41][29] = -8'd7;
        rom[41][30] = -8'd3;
        rom[41][31] = 8'd9;
        rom[42][0] = -8'd30;
        rom[42][1] = 8'd16;
        rom[42][2] = 8'd9;
        rom[42][3] = 8'd23;
        rom[42][4] = -8'd11;
        rom[42][5] = -8'd37;
        rom[42][6] = -8'd14;
        rom[42][7] = 8'd4;
        rom[42][8] = 8'd14;
        rom[42][9] = -8'd19;
        rom[42][10] = 8'd31;
        rom[42][11] = 8'd16;
        rom[42][12] = -8'd18;
        rom[42][13] = 8'd19;
        rom[42][14] = -8'd9;
        rom[42][15] = -8'd20;
        rom[42][16] = -8'd2;
        rom[42][17] = -8'd47;
        rom[42][18] = 8'd13;
        rom[42][19] = 8'd3;
        rom[42][20] = -8'd6;
        rom[42][21] = -8'd6;
        rom[42][22] = 8'd0;
        rom[42][23] = 8'd12;
        rom[42][24] = 8'd26;
        rom[42][25] = -8'd21;
        rom[42][26] = 8'd54;
        rom[42][27] = -8'd15;
        rom[42][28] = 8'd23;
        rom[42][29] = -8'd5;
        rom[42][30] = 8'd9;
        rom[42][31] = -8'd26;
        rom[43][0] = 8'd8;
        rom[43][1] = 8'd3;
        rom[43][2] = -8'd30;
        rom[43][3] = 8'd49;
        rom[43][4] = 8'd13;
        rom[43][5] = -8'd23;
        rom[43][6] = 8'd1;
        rom[43][7] = -8'd20;
        rom[43][8] = -8'd5;
        rom[43][9] = -8'd2;
        rom[43][10] = -8'd6;
        rom[43][11] = 8'd10;
        rom[43][12] = 8'd24;
        rom[43][13] = 8'd26;
        rom[43][14] = 8'd32;
        rom[43][15] = 8'd20;
        rom[43][16] = 8'd2;
        rom[43][17] = -8'd9;
        rom[43][18] = -8'd39;
        rom[43][19] = 8'd4;
        rom[43][20] = -8'd27;
        rom[43][21] = 8'd24;
        rom[43][22] = -8'd26;
        rom[43][23] = -8'd6;
        rom[43][24] = -8'd1;
        rom[43][25] = 8'd3;
        rom[43][26] = -8'd1;
        rom[43][27] = -8'd24;
        rom[43][28] = 8'd7;
        rom[43][29] = -8'd38;
        rom[43][30] = -8'd6;
        rom[43][31] = 8'd38;
        rom[44][0] = 8'd20;
        rom[44][1] = -8'd19;
        rom[44][2] = 8'd21;
        rom[44][3] = -8'd20;
        rom[44][4] = 8'd28;
        rom[44][5] = -8'd2;
        rom[44][6] = 8'd27;
        rom[44][7] = 8'd19;
        rom[44][8] = -8'd1;
        rom[44][9] = 8'd25;
        rom[44][10] = 8'd9;
        rom[44][11] = 8'd12;
        rom[44][12] = 8'd6;
        rom[44][13] = -8'd58;
        rom[44][14] = 8'd9;
        rom[44][15] = -8'd8;
        rom[44][16] = 8'd7;
        rom[44][17] = 8'd9;
        rom[44][18] = -8'd35;
        rom[44][19] = 8'd33;
        rom[44][20] = -8'd10;
        rom[44][21] = 8'd19;
        rom[44][22] = -8'd60;
        rom[44][23] = 8'd2;
        rom[44][24] = -8'd15;
        rom[44][25] = 8'd16;
        rom[44][26] = 8'd18;
        rom[44][27] = 8'd13;
        rom[44][28] = -8'd6;
        rom[44][29] = 8'd37;
        rom[44][30] = 8'd3;
        rom[44][31] = 8'd15;
        rom[45][0] = 8'd0;
        rom[45][1] = 8'd13;
        rom[45][2] = -8'd7;
        rom[45][3] = 8'd14;
        rom[45][4] = 8'd20;
        rom[45][5] = -8'd8;
        rom[45][6] = 8'd0;
        rom[45][7] = -8'd7;
        rom[45][8] = 8'd19;
        rom[45][9] = -8'd18;
        rom[45][10] = -8'd6;
        rom[45][11] = -8'd4;
        rom[45][12] = -8'd37;
        rom[45][13] = -8'd24;
        rom[45][14] = -8'd35;
        rom[45][15] = 8'd19;
        rom[45][16] = -8'd18;
        rom[45][17] = -8'd18;
        rom[45][18] = -8'd3;
        rom[45][19] = 8'd5;
        rom[45][20] = 8'd15;
        rom[45][21] = -8'd19;
        rom[45][22] = 8'd8;
        rom[45][23] = -8'd9;
        rom[45][24] = 8'd23;
        rom[45][25] = -8'd16;
        rom[45][26] = 8'd17;
        rom[45][27] = 8'd23;
        rom[45][28] = -8'd29;
        rom[45][29] = 8'd16;
        rom[45][30] = 8'd13;
        rom[45][31] = 8'd22;
        rom[46][0] = 8'd16;
        rom[46][1] = 8'd34;
        rom[46][2] = 8'd18;
        rom[46][3] = 8'd1;
        rom[46][4] = -8'd42;
        rom[46][5] = -8'd17;
        rom[46][6] = -8'd1;
        rom[46][7] = 8'd6;
        rom[46][8] = -8'd19;
        rom[46][9] = -8'd21;
        rom[46][10] = 8'd20;
        rom[46][11] = -8'd24;
        rom[46][12] = 8'd29;
        rom[46][13] = -8'd41;
        rom[46][14] = -8'd11;
        rom[46][15] = -8'd8;
        rom[46][16] = 8'd16;
        rom[46][17] = -8'd4;
        rom[46][18] = 8'd30;
        rom[46][19] = 8'd30;
        rom[46][20] = 8'd31;
        rom[46][21] = 8'd6;
        rom[46][22] = -8'd51;
        rom[46][23] = 8'd30;
        rom[46][24] = 8'd11;
        rom[46][25] = -8'd32;
        rom[46][26] = -8'd26;
        rom[46][27] = 8'd9;
        rom[46][28] = -8'd3;
        rom[46][29] = -8'd32;
        rom[46][30] = -8'd13;
        rom[46][31] = 8'd34;
        rom[47][0] = -8'd19;
        rom[47][1] = -8'd20;
        rom[47][2] = -8'd19;
        rom[47][3] = 8'd13;
        rom[47][4] = 8'd9;
        rom[47][5] = -8'd53;
        rom[47][6] = 8'd19;
        rom[47][7] = 8'd4;
        rom[47][8] = -8'd4;
        rom[47][9] = -8'd26;
        rom[47][10] = -8'd24;
        rom[47][11] = -8'd4;
        rom[47][12] = 8'd27;
        rom[47][13] = -8'd20;
        rom[47][14] = 8'd9;
        rom[47][15] = -8'd15;
        rom[47][16] = 8'd12;
        rom[47][17] = -8'd35;
        rom[47][18] = 8'd2;
        rom[47][19] = 8'd0;
        rom[47][20] = 8'd28;
        rom[47][21] = -8'd16;
        rom[47][22] = -8'd14;
        rom[47][23] = 8'd12;
        rom[47][24] = 8'd26;
        rom[47][25] = 8'd21;
        rom[47][26] = 8'd23;
        rom[47][27] = -8'd7;
        rom[47][28] = 8'd22;
        rom[47][29] = -8'd4;
        rom[47][30] = 8'd7;
        rom[47][31] = 8'd0;
        rom[48][0] = -8'd19;
        rom[48][1] = 8'd4;
        rom[48][2] = 8'd11;
        rom[48][3] = -8'd36;
        rom[48][4] = 8'd19;
        rom[48][5] = 8'd0;
        rom[48][6] = -8'd3;
        rom[48][7] = 8'd18;
        rom[48][8] = 8'd16;
        rom[48][9] = 8'd12;
        rom[48][10] = -8'd30;
        rom[48][11] = -8'd51;
        rom[48][12] = 8'd11;
        rom[48][13] = 8'd0;
        rom[48][14] = 8'd12;
        rom[48][15] = -8'd22;
        rom[48][16] = -8'd9;
        rom[48][17] = -8'd1;
        rom[48][18] = 8'd23;
        rom[48][19] = 8'd8;
        rom[48][20] = 8'd2;
        rom[48][21] = 8'd3;
        rom[48][22] = 8'd13;
        rom[48][23] = -8'd30;
        rom[48][24] = -8'd19;
        rom[48][25] = 8'd24;
        rom[48][26] = -8'd12;
        rom[48][27] = -8'd17;
        rom[48][28] = 8'd9;
        rom[48][29] = 8'd36;
        rom[48][30] = -8'd17;
        rom[48][31] = -8'd18;
        rom[49][0] = -8'd9;
        rom[49][1] = -8'd15;
        rom[49][2] = -8'd11;
        rom[49][3] = 8'd14;
        rom[49][4] = 8'd28;
        rom[49][5] = -8'd9;
        rom[49][6] = -8'd2;
        rom[49][7] = -8'd8;
        rom[49][8] = 8'd27;
        rom[49][9] = -8'd35;
        rom[49][10] = -8'd21;
        rom[49][11] = -8'd14;
        rom[49][12] = 8'd1;
        rom[49][13] = 8'd3;
        rom[49][14] = -8'd24;
        rom[49][15] = 8'd12;
        rom[49][16] = 8'd7;
        rom[49][17] = -8'd33;
        rom[49][18] = 8'd3;
        rom[49][19] = 8'd13;
        rom[49][20] = -8'd48;
        rom[49][21] = 8'd3;
        rom[49][22] = -8'd9;
        rom[49][23] = -8'd8;
        rom[49][24] = 8'd10;
        rom[49][25] = 8'd17;
        rom[49][26] = 8'd12;
        rom[49][27] = -8'd37;
        rom[49][28] = -8'd46;
        rom[49][29] = -8'd36;
        rom[49][30] = -8'd15;
        rom[49][31] = -8'd11;
        rom[50][0] = 8'd14;
        rom[50][1] = 8'd46;
        rom[50][2] = -8'd1;
        rom[50][3] = -8'd21;
        rom[50][4] = -8'd11;
        rom[50][5] = 8'd0;
        rom[50][6] = 8'd2;
        rom[50][7] = -8'd14;
        rom[50][8] = 8'd34;
        rom[50][9] = -8'd5;
        rom[50][10] = -8'd17;
        rom[50][11] = -8'd22;
        rom[50][12] = 8'd4;
        rom[50][13] = -8'd7;
        rom[50][14] = 8'd19;
        rom[50][15] = 8'd6;
        rom[50][16] = 8'd4;
        rom[50][17] = 8'd7;
        rom[50][18] = -8'd11;
        rom[50][19] = 8'd8;
        rom[50][20] = -8'd13;
        rom[50][21] = -8'd20;
        rom[50][22] = -8'd6;
        rom[50][23] = 8'd27;
        rom[50][24] = 8'd0;
        rom[50][25] = 8'd17;
        rom[50][26] = 8'd5;
        rom[50][27] = -8'd15;
        rom[50][28] = -8'd25;
        rom[50][29] = -8'd17;
        rom[50][30] = -8'd34;
        rom[50][31] = 8'd2;
        rom[51][0] = 8'd12;
        rom[51][1] = 8'd62;
        rom[51][2] = 8'd17;
        rom[51][3] = -8'd14;
        rom[51][4] = 8'd44;
        rom[51][5] = -8'd9;
        rom[51][6] = -8'd12;
        rom[51][7] = -8'd5;
        rom[51][8] = 8'd44;
        rom[51][9] = -8'd8;
        rom[51][10] = -8'd36;
        rom[51][11] = -8'd23;
        rom[51][12] = -8'd11;
        rom[51][13] = -8'd5;
        rom[51][14] = -8'd6;
        rom[51][15] = 8'd10;
        rom[51][16] = 8'd3;
        rom[51][17] = -8'd12;
        rom[51][18] = 8'd27;
        rom[51][19] = 8'd10;
        rom[51][20] = -8'd24;
        rom[51][21] = -8'd13;
        rom[51][22] = 8'd4;
        rom[51][23] = 8'd21;
        rom[51][24] = 8'd10;
        rom[51][25] = 8'd25;
        rom[51][26] = -8'd36;
        rom[51][27] = 8'd10;
        rom[51][28] = -8'd19;
        rom[51][29] = 8'd13;
        rom[51][30] = -8'd44;
        rom[51][31] = 8'd15;
        rom[52][0] = 8'd29;
        rom[52][1] = 8'd35;
        rom[52][2] = 8'd1;
        rom[52][3] = -8'd5;
        rom[52][4] = 8'd38;
        rom[52][5] = -8'd24;
        rom[52][6] = -8'd39;
        rom[52][7] = 8'd14;
        rom[52][8] = 8'd48;
        rom[52][9] = -8'd7;
        rom[52][10] = 8'd9;
        rom[52][11] = -8'd109;
        rom[52][12] = 8'd7;
        rom[52][13] = 8'd19;
        rom[52][14] = -8'd4;
        rom[52][15] = 8'd20;
        rom[52][16] = -8'd5;
        rom[52][17] = 8'd1;
        rom[52][18] = 8'd21;
        rom[52][19] = 8'd3;
        rom[52][20] = -8'd33;
        rom[52][21] = 8'd11;
        rom[52][22] = 8'd26;
        rom[52][23] = -8'd41;
        rom[52][24] = -8'd21;
        rom[52][25] = 8'd30;
        rom[52][26] = 8'd18;
        rom[52][27] = 8'd5;
        rom[52][28] = -8'd3;
        rom[52][29] = -8'd73;
        rom[52][30] = -8'd3;
        rom[52][31] = 8'd10;
        rom[53][0] = -8'd24;
        rom[53][1] = 8'd9;
        rom[53][2] = -8'd16;
        rom[53][3] = 8'd23;
        rom[53][4] = -8'd15;
        rom[53][5] = 8'd23;
        rom[53][6] = 8'd21;
        rom[53][7] = 8'd21;
        rom[53][8] = 8'd27;
        rom[53][9] = -8'd16;
        rom[53][10] = -8'd67;
        rom[53][11] = 8'd1;
        rom[53][12] = -8'd5;
        rom[53][13] = -8'd22;
        rom[53][14] = 8'd20;
        rom[53][15] = -8'd13;
        rom[53][16] = 8'd18;
        rom[53][17] = 8'd2;
        rom[53][18] = -8'd57;
        rom[53][19] = -8'd33;
        rom[53][20] = 8'd17;
        rom[53][21] = 8'd27;
        rom[53][22] = 8'd20;
        rom[53][23] = 8'd13;
        rom[53][24] = -8'd12;
        rom[53][25] = 8'd11;
        rom[53][26] = 8'd14;
        rom[53][27] = -8'd1;
        rom[53][28] = 8'd15;
        rom[53][29] = 8'd15;
        rom[53][30] = 8'd5;
        rom[53][31] = -8'd59;
        rom[54][0] = 8'd13;
        rom[54][1] = 8'd24;
        rom[54][2] = 8'd0;
        rom[54][3] = -8'd16;
        rom[54][4] = -8'd12;
        rom[54][5] = -8'd21;
        rom[54][6] = 8'd1;
        rom[54][7] = 8'd1;
        rom[54][8] = 8'd6;
        rom[54][9] = 8'd14;
        rom[54][10] = 8'd12;
        rom[54][11] = -8'd52;
        rom[54][12] = -8'd1;
        rom[54][13] = 8'd13;
        rom[54][14] = 8'd0;
        rom[54][15] = 8'd31;
        rom[54][16] = -8'd50;
        rom[54][17] = -8'd19;
        rom[54][18] = -8'd6;
        rom[54][19] = -8'd9;
        rom[54][20] = -8'd4;
        rom[54][21] = -8'd40;
        rom[54][22] = -8'd33;
        rom[54][23] = 8'd21;
        rom[54][24] = -8'd28;
        rom[54][25] = 8'd4;
        rom[54][26] = -8'd5;
        rom[54][27] = 8'd22;
        rom[54][28] = 8'd14;
        rom[54][29] = 8'd5;
        rom[54][30] = 8'd9;
        rom[54][31] = 8'd24;
        rom[55][0] = 8'd0;
        rom[55][1] = 8'd0;
        rom[55][2] = 8'd1;
        rom[55][3] = -8'd18;
        rom[55][4] = 8'd4;
        rom[55][5] = 8'd20;
        rom[55][6] = -8'd13;
        rom[55][7] = -8'd17;
        rom[55][8] = 8'd23;
        rom[55][9] = -8'd60;
        rom[55][10] = 8'd7;
        rom[55][11] = -8'd7;
        rom[55][12] = 8'd8;
        rom[55][13] = -8'd14;
        rom[55][14] = -8'd23;
        rom[55][15] = -8'd46;
        rom[55][16] = 8'd1;
        rom[55][17] = -8'd7;
        rom[55][18] = -8'd10;
        rom[55][19] = 8'd10;
        rom[55][20] = 8'd20;
        rom[55][21] = -8'd6;
        rom[55][22] = -8'd1;
        rom[55][23] = 8'd1;
        rom[55][24] = 8'd2;
        rom[55][25] = 8'd2;
        rom[55][26] = 8'd3;
        rom[55][27] = 8'd16;
        rom[55][28] = 8'd13;
        rom[55][29] = 8'd1;
        rom[55][30] = 8'd16;
        rom[55][31] = -8'd45;
        rom[56][0] = 8'd17;
        rom[56][1] = 8'd22;
        rom[56][2] = 8'd39;
        rom[56][3] = -8'd15;
        rom[56][4] = -8'd7;
        rom[56][5] = -8'd16;
        rom[56][6] = 8'd12;
        rom[56][7] = -8'd6;
        rom[56][8] = 8'd34;
        rom[56][9] = -8'd6;
        rom[56][10] = 8'd6;
        rom[56][11] = -8'd58;
        rom[56][12] = 8'd10;
        rom[56][13] = -8'd5;
        rom[56][14] = 8'd5;
        rom[56][15] = 8'd1;
        rom[56][16] = -8'd34;
        rom[56][17] = -8'd12;
        rom[56][18] = 8'd16;
        rom[56][19] = -8'd67;
        rom[56][20] = -8'd7;
        rom[56][21] = -8'd10;
        rom[56][22] = -8'd24;
        rom[56][23] = -8'd14;
        rom[56][24] = -8'd41;
        rom[56][25] = -8'd12;
        rom[56][26] = 8'd2;
        rom[56][27] = -8'd8;
        rom[56][28] = 8'd24;
        rom[56][29] = -8'd3;
        rom[56][30] = -8'd16;
        rom[56][31] = 8'd3;
        rom[57][0] = -8'd4;
        rom[57][1] = -8'd39;
        rom[57][2] = 8'd44;
        rom[57][3] = -8'd25;
        rom[57][4] = -8'd33;
        rom[57][5] = 8'd10;
        rom[57][6] = 8'd13;
        rom[57][7] = 8'd33;
        rom[57][8] = -8'd21;
        rom[57][9] = 8'd27;
        rom[57][10] = -8'd3;
        rom[57][11] = -8'd37;
        rom[57][12] = 8'd4;
        rom[57][13] = 8'd11;
        rom[57][14] = 8'd0;
        rom[57][15] = 8'd17;
        rom[57][16] = 8'd16;
        rom[57][17] = 8'd19;
        rom[57][18] = 8'd16;
        rom[57][19] = -8'd25;
        rom[57][20] = -8'd8;
        rom[57][21] = -8'd57;
        rom[57][22] = 8'd15;
        rom[57][23] = -8'd10;
        rom[57][24] = -8'd17;
        rom[57][25] = -8'd3;
        rom[57][26] = 8'd10;
        rom[57][27] = 8'd23;
        rom[57][28] = -8'd23;
        rom[57][29] = 8'd7;
        rom[57][30] = 8'd40;
        rom[57][31] = -8'd1;
        rom[58][0] = -8'd6;
        rom[58][1] = 8'd51;
        rom[58][2] = -8'd9;
        rom[58][3] = 8'd29;
        rom[58][4] = 8'd0;
        rom[58][5] = -8'd35;
        rom[58][6] = 8'd6;
        rom[58][7] = -8'd4;
        rom[58][8] = 8'd11;
        rom[58][9] = 8'd8;
        rom[58][10] = 8'd1;
        rom[58][11] = 8'd1;
        rom[58][12] = 8'd19;
        rom[58][13] = 8'd43;
        rom[58][14] = 8'd22;
        rom[58][15] = 8'd24;
        rom[58][16] = -8'd23;
        rom[58][17] = -8'd8;
        rom[58][18] = 8'd28;
        rom[58][19] = 8'd49;
        rom[58][20] = -8'd79;
        rom[58][21] = -8'd51;
        rom[58][22] = 8'd39;
        rom[58][23] = 8'd29;
        rom[58][24] = -8'd31;
        rom[58][25] = 8'd33;
        rom[58][26] = 8'd24;
        rom[58][27] = 8'd11;
        rom[58][28] = 8'd18;
        rom[58][29] = -8'd17;
        rom[58][30] = -8'd50;
        rom[58][31] = 8'd6;
        rom[59][0] = -8'd38;
        rom[59][1] = -8'd10;
        rom[59][2] = 8'd10;
        rom[59][3] = -8'd17;
        rom[59][4] = -8'd1;
        rom[59][5] = 8'd10;
        rom[59][6] = 8'd4;
        rom[59][7] = 8'd25;
        rom[59][8] = 8'd3;
        rom[59][9] = -8'd2;
        rom[59][10] = -8'd60;
        rom[59][11] = 8'd27;
        rom[59][12] = -8'd13;
        rom[59][13] = 8'd0;
        rom[59][14] = 8'd12;
        rom[59][15] = 8'd4;
        rom[59][16] = -8'd13;
        rom[59][17] = -8'd38;
        rom[59][18] = -8'd44;
        rom[59][19] = -8'd11;
        rom[59][20] = -8'd3;
        rom[59][21] = 8'd23;
        rom[59][22] = 8'd16;
        rom[59][23] = 8'd10;
        rom[59][24] = -8'd4;
        rom[59][25] = 8'd29;
        rom[59][26] = 8'd0;
        rom[59][27] = 8'd15;
        rom[59][28] = 8'd20;
        rom[59][29] = 8'd0;
        rom[59][30] = 8'd5;
        rom[59][31] = -8'd30;
        rom[60][0] = 8'd9;
        rom[60][1] = -8'd2;
        rom[60][2] = 8'd10;
        rom[60][3] = 8'd41;
        rom[60][4] = -8'd17;
        rom[60][5] = 8'd3;
        rom[60][6] = -8'd31;
        rom[60][7] = 8'd14;
        rom[60][8] = 8'd25;
        rom[60][9] = 8'd11;
        rom[60][10] = -8'd20;
        rom[60][11] = -8'd29;
        rom[60][12] = 8'd7;
        rom[60][13] = -8'd22;
        rom[60][14] = 8'd1;
        rom[60][15] = 8'd27;
        rom[60][16] = 8'd21;
        rom[60][17] = -8'd5;
        rom[60][18] = -8'd18;
        rom[60][19] = -8'd9;
        rom[60][20] = 8'd32;
        rom[60][21] = -8'd34;
        rom[60][22] = -8'd38;
        rom[60][23] = -8'd17;
        rom[60][24] = 8'd23;
        rom[60][25] = -8'd8;
        rom[60][26] = -8'd12;
        rom[60][27] = -8'd15;
        rom[60][28] = -8'd11;
        rom[60][29] = 8'd12;
        rom[60][30] = 8'd44;
        rom[60][31] = -8'd20;
        rom[61][0] = -8'd5;
        rom[61][1] = -8'd11;
        rom[61][2] = 8'd5;
        rom[61][3] = 8'd0;
        rom[61][4] = -8'd33;
        rom[61][5] = 8'd1;
        rom[61][6] = 8'd0;
        rom[61][7] = 8'd15;
        rom[61][8] = 8'd4;
        rom[61][9] = 8'd40;
        rom[61][10] = -8'd72;
        rom[61][11] = -8'd7;
        rom[61][12] = 8'd21;
        rom[61][13] = -8'd33;
        rom[61][14] = 8'd5;
        rom[61][15] = 8'd0;
        rom[61][16] = -8'd15;
        rom[61][17] = 8'd8;
        rom[61][18] = -8'd32;
        rom[61][19] = -8'd14;
        rom[61][20] = 8'd2;
        rom[61][21] = 8'd14;
        rom[61][22] = -8'd9;
        rom[61][23] = 8'd17;
        rom[61][24] = -8'd22;
        rom[61][25] = -8'd17;
        rom[61][26] = -8'd21;
        rom[61][27] = 8'd21;
        rom[61][28] = 8'd2;
        rom[61][29] = 8'd20;
        rom[61][30] = 8'd12;
        rom[61][31] = -8'd17;
        rom[62][0] = -8'd26;
        rom[62][1] = -8'd13;
        rom[62][2] = 8'd6;
        rom[62][3] = 8'd11;
        rom[62][4] = -8'd4;
        rom[62][5] = 8'd6;
        rom[62][6] = 8'd15;
        rom[62][7] = 8'd4;
        rom[62][8] = 8'd16;
        rom[62][9] = 8'd3;
        rom[62][10] = -8'd14;
        rom[62][11] = 8'd12;
        rom[62][12] = 8'd20;
        rom[62][13] = 8'd23;
        rom[62][14] = -8'd6;
        rom[62][15] = -8'd22;
        rom[62][16] = -8'd45;
        rom[62][17] = 8'd10;
        rom[62][18] = -8'd9;
        rom[62][19] = 8'd21;
        rom[62][20] = -8'd21;
        rom[62][21] = -8'd6;
        rom[62][22] = 8'd14;
        rom[62][23] = -8'd13;
        rom[62][24] = 8'd8;
        rom[62][25] = 8'd28;
        rom[62][26] = 8'd22;
        rom[62][27] = -8'd14;
        rom[62][28] = 8'd23;
        rom[62][29] = 8'd8;
        rom[62][30] = 8'd16;
        rom[62][31] = -8'd5;
        rom[63][0] = -8'd23;
        rom[63][1] = 8'd38;
        rom[63][2] = -8'd52;
        rom[63][3] = 8'd15;
        rom[63][4] = -8'd30;
        rom[63][5] = 8'd19;
        rom[63][6] = 8'd5;
        rom[63][7] = 8'd1;
        rom[63][8] = 8'd18;
        rom[63][9] = 8'd22;
        rom[63][10] = -8'd19;
        rom[63][11] = -8'd24;
        rom[63][12] = 8'd7;
        rom[63][13] = -8'd22;
        rom[63][14] = -8'd2;
        rom[63][15] = 8'd14;
        rom[63][16] = -8'd14;
        rom[63][17] = 8'd28;
        rom[63][18] = -8'd72;
        rom[63][19] = 8'd6;
        rom[63][20] = -8'd2;
        rom[63][21] = 8'd24;
        rom[63][22] = -8'd4;
        rom[63][23] = 8'd14;
        rom[63][24] = 8'd14;
        rom[63][25] = 8'd5;
        rom[63][26] = 8'd7;
        rom[63][27] = 8'd30;
        rom[63][28] = -8'd13;
        rom[63][29] = 8'd26;
        rom[63][30] = -8'd28;
        rom[63][31] = -8'd16;
        rom[64][0] = 8'd1;
        rom[64][1] = -8'd45;
        rom[64][2] = 8'd18;
        rom[64][3] = -8'd76;
        rom[64][4] = 8'd26;
        rom[64][5] = -8'd29;
        rom[64][6] = -8'd27;
        rom[64][7] = 8'd1;
        rom[64][8] = 8'd13;
        rom[64][9] = 8'd0;
        rom[64][10] = 8'd10;
        rom[64][11] = -8'd32;
        rom[64][12] = 8'd0;
        rom[64][13] = 8'd0;
        rom[64][14] = -8'd6;
        rom[64][15] = 8'd26;
        rom[64][16] = -8'd14;
        rom[64][17] = 8'd42;
        rom[64][18] = 8'd7;
        rom[64][19] = -8'd20;
        rom[64][20] = -8'd13;
        rom[64][21] = -8'd14;
        rom[64][22] = 8'd5;
        rom[64][23] = -8'd4;
        rom[64][24] = -8'd97;
        rom[64][25] = -8'd5;
        rom[64][26] = 8'd1;
        rom[64][27] = -8'd59;
        rom[64][28] = 8'd24;
        rom[64][29] = 8'd10;
        rom[64][30] = -8'd32;
        rom[64][31] = -8'd17;
        rom[65][0] = 8'd4;
        rom[65][1] = 8'd0;
        rom[65][2] = -8'd23;
        rom[65][3] = 8'd48;
        rom[65][4] = 8'd5;
        rom[65][5] = 8'd5;
        rom[65][6] = -8'd4;
        rom[65][7] = 8'd0;
        rom[65][8] = -8'd2;
        rom[65][9] = 8'd0;
        rom[65][10] = 8'd14;
        rom[65][11] = -8'd11;
        rom[65][12] = 8'd41;
        rom[65][13] = 8'd24;
        rom[65][14] = -8'd20;
        rom[65][15] = 8'd18;
        rom[65][16] = 8'd43;
        rom[65][17] = -8'd34;
        rom[65][18] = 8'd9;
        rom[65][19] = 8'd18;
        rom[65][20] = -8'd22;
        rom[65][21] = 8'd23;
        rom[65][22] = -8'd36;
        rom[65][23] = -8'd7;
        rom[65][24] = 8'd7;
        rom[65][25] = 8'd17;
        rom[65][26] = 8'd0;
        rom[65][27] = -8'd8;
        rom[65][28] = 8'd7;
        rom[65][29] = -8'd14;
        rom[65][30] = 8'd12;
        rom[65][31] = -8'd31;
        rom[66][0] = -8'd8;
        rom[66][1] = 8'd29;
        rom[66][2] = -8'd47;
        rom[66][3] = 8'd0;
        rom[66][4] = 8'd5;
        rom[66][5] = -8'd17;
        rom[66][6] = -8'd27;
        rom[66][7] = 8'd22;
        rom[66][8] = 8'd30;
        rom[66][9] = -8'd45;
        rom[66][10] = -8'd26;
        rom[66][11] = 8'd22;
        rom[66][12] = -8'd29;
        rom[66][13] = 8'd15;
        rom[66][14] = 8'd9;
        rom[66][15] = -8'd12;
        rom[66][16] = 8'd35;
        rom[66][17] = -8'd68;
        rom[66][18] = -8'd3;
        rom[66][19] = 8'd37;
        rom[66][20] = -8'd6;
        rom[66][21] = -8'd19;
        rom[66][22] = 8'd10;
        rom[66][23] = 8'd32;
        rom[66][24] = -8'd4;
        rom[66][25] = 8'd4;
        rom[66][26] = -8'd17;
        rom[66][27] = 8'd13;
        rom[66][28] = -8'd40;
        rom[66][29] = 8'd11;
        rom[66][30] = -8'd45;
        rom[66][31] = 8'd15;
        rom[67][0] = 8'd25;
        rom[67][1] = -8'd11;
        rom[67][2] = 8'd27;
        rom[67][3] = -8'd7;
        rom[67][4] = 8'd27;
        rom[67][5] = 8'd31;
        rom[67][6] = -8'd29;
        rom[67][7] = -8'd1;
        rom[67][8] = 8'd18;
        rom[67][9] = 8'd20;
        rom[67][10] = -8'd4;
        rom[67][11] = -8'd12;
        rom[67][12] = 8'd48;
        rom[67][13] = 8'd2;
        rom[67][14] = -8'd22;
        rom[67][15] = 8'd8;
        rom[67][16] = 8'd29;
        rom[67][17] = 8'd4;
        rom[67][18] = 8'd24;
        rom[67][19] = -8'd20;
        rom[67][20] = 8'd17;
        rom[67][21] = -8'd26;
        rom[67][22] = 8'd26;
        rom[67][23] = -8'd43;
        rom[67][24] = 8'd13;
        rom[67][25] = 8'd32;
        rom[67][26] = -8'd55;
        rom[67][27] = -8'd8;
        rom[67][28] = 8'd19;
        rom[67][29] = -8'd32;
        rom[67][30] = 8'd33;
        rom[67][31] = -8'd1;
        rom[68][0] = 8'd32;
        rom[68][1] = -8'd45;
        rom[68][2] = 8'd7;
        rom[68][3] = -8'd1;
        rom[68][4] = 8'd46;
        rom[68][5] = -8'd3;
        rom[68][6] = -8'd84;
        rom[68][7] = 8'd13;
        rom[68][8] = 8'd34;
        rom[68][9] = 8'd5;
        rom[68][10] = -8'd10;
        rom[68][11] = -8'd18;
        rom[68][12] = -8'd4;
        rom[68][13] = 8'd7;
        rom[68][14] = -8'd16;
        rom[68][15] = 8'd31;
        rom[68][16] = 8'd13;
        rom[68][17] = 8'd36;
        rom[68][18] = 8'd23;
        rom[68][19] = -8'd31;
        rom[68][20] = -8'd24;
        rom[68][21] = -8'd10;
        rom[68][22] = 8'd31;
        rom[68][23] = -8'd17;
        rom[68][24] = -8'd116;
        rom[68][25] = 8'd2;
        rom[68][26] = 8'd18;
        rom[68][27] = -8'd11;
        rom[68][28] = 8'd9;
        rom[68][29] = -8'd75;
        rom[68][30] = 8'd39;
        rom[68][31] = 8'd18;
        rom[69][0] = -8'd9;
        rom[69][1] = 8'd15;
        rom[69][2] = -8'd112;
        rom[69][3] = -8'd32;
        rom[69][4] = -8'd5;
        rom[69][5] = 8'd12;
        rom[69][6] = 8'd14;
        rom[69][7] = 8'd26;
        rom[69][8] = 8'd1;
        rom[69][9] = -8'd110;
        rom[69][10] = -8'd15;
        rom[69][11] = 8'd29;
        rom[69][12] = -8'd55;
        rom[69][13] = -8'd64;
        rom[69][14] = -8'd12;
        rom[69][15] = -8'd19;
        rom[69][16] = 8'd16;
        rom[69][17] = 8'd13;
        rom[69][18] = -8'd94;
        rom[69][19] = -8'd85;
        rom[69][20] = 8'd6;
        rom[69][21] = 8'd22;
        rom[69][22] = 8'd13;
        rom[69][23] = 8'd25;
        rom[69][24] = -8'd1;
        rom[69][25] = 8'd17;
        rom[69][26] = 8'd7;
        rom[69][27] = 8'd0;
        rom[69][28] = -8'd51;
        rom[69][29] = 8'd31;
        rom[69][30] = 8'd15;
        rom[69][31] = -8'd58;
        rom[70][0] = 8'd1;
        rom[70][1] = -8'd48;
        rom[70][2] = -8'd29;
        rom[70][3] = 8'd27;
        rom[70][4] = 8'd8;
        rom[70][5] = -8'd78;
        rom[70][6] = -8'd56;
        rom[70][7] = 8'd21;
        rom[70][8] = 8'd3;
        rom[70][9] = 8'd27;
        rom[70][10] = -8'd29;
        rom[70][11] = -8'd9;
        rom[70][12] = 8'd5;
        rom[70][13] = 8'd13;
        rom[70][14] = 8'd27;
        rom[70][15] = 8'd9;
        rom[70][16] = -8'd41;
        rom[70][17] = -8'd8;
        rom[70][18] = -8'd4;
        rom[70][19] = 8'd40;
        rom[70][20] = -8'd4;
        rom[70][21] = -8'd10;
        rom[70][22] = -8'd25;
        rom[70][23] = -8'd2;
        rom[70][24] = -8'd128;
        rom[70][25] = -8'd78;
        rom[70][26] = -8'd28;
        rom[70][27] = 8'd23;
        rom[70][28] = 8'd7;
        rom[70][29] = -8'd10;
        rom[70][30] = 8'd37;
        rom[70][31] = 8'd21;
        rom[71][0] = -8'd29;
        rom[71][1] = -8'd12;
        rom[71][2] = -8'd6;
        rom[71][3] = -8'd57;
        rom[71][4] = -8'd31;
        rom[71][5] = 8'd10;
        rom[71][6] = 8'd16;
        rom[71][7] = 8'd36;
        rom[71][8] = -8'd8;
        rom[71][9] = -8'd33;
        rom[71][10] = 8'd40;
        rom[71][11] = 8'd25;
        rom[71][12] = -8'd15;
        rom[71][13] = -8'd41;
        rom[71][14] = -8'd32;
        rom[71][15] = -8'd34;
        rom[71][16] = -8'd12;
        rom[71][17] = 8'd47;
        rom[71][18] = -8'd46;
        rom[71][19] = -8'd17;
        rom[71][20] = 8'd22;
        rom[71][21] = 8'd11;
        rom[71][22] = 8'd6;
        rom[71][23] = 8'd21;
        rom[71][24] = 8'd9;
        rom[71][25] = 8'd32;
        rom[71][26] = -8'd22;
        rom[71][27] = 8'd14;
        rom[71][28] = -8'd23;
        rom[71][29] = 8'd7;
        rom[71][30] = 8'd20;
        rom[71][31] = -8'd34;
        rom[72][0] = 8'd34;
        rom[72][1] = -8'd31;
        rom[72][2] = 8'd30;
        rom[72][3] = -8'd3;
        rom[72][4] = -8'd18;
        rom[72][5] = -8'd48;
        rom[72][6] = 8'd22;
        rom[72][7] = 8'd36;
        rom[72][8] = 8'd1;
        rom[72][9] = 8'd7;
        rom[72][10] = 8'd6;
        rom[72][11] = -8'd21;
        rom[72][12] = -8'd20;
        rom[72][13] = 8'd19;
        rom[72][14] = 8'd12;
        rom[72][15] = 8'd15;
        rom[72][16] = -8'd35;
        rom[72][17] = 8'd38;
        rom[72][18] = 8'd19;
        rom[72][19] = -8'd103;
        rom[72][20] = -8'd20;
        rom[72][21] = -8'd19;
        rom[72][22] = -8'd14;
        rom[72][23] = 8'd21;
        rom[72][24] = -8'd128;
        rom[72][25] = -8'd21;
        rom[72][26] = 8'd9;
        rom[72][27] = -8'd10;
        rom[72][28] = 8'd28;
        rom[72][29] = -8'd18;
        rom[72][30] = 8'd7;
        rom[72][31] = -8'd4;
        rom[73][0] = -8'd6;
        rom[73][1] = -8'd60;
        rom[73][2] = 8'd2;
        rom[73][3] = 8'd12;
        rom[73][4] = -8'd20;
        rom[73][5] = -8'd19;
        rom[73][6] = 8'd43;
        rom[73][7] = 8'd4;
        rom[73][8] = -8'd31;
        rom[73][9] = -8'd19;
        rom[73][10] = 8'd4;
        rom[73][11] = -8'd50;
        rom[73][12] = 8'd27;
        rom[73][13] = -8'd38;
        rom[73][14] = -8'd31;
        rom[73][15] = 8'd54;
        rom[73][16] = 8'd9;
        rom[73][17] = 8'd21;
        rom[73][18] = 8'd10;
        rom[73][19] = -8'd32;
        rom[73][20] = -8'd42;
        rom[73][21] = -8'd74;
        rom[73][22] = 8'd27;
        rom[73][23] = -8'd26;
        rom[73][24] = -8'd85;
        rom[73][25] = 8'd6;
        rom[73][26] = 8'd18;
        rom[73][27] = -8'd3;
        rom[73][28] = -8'd20;
        rom[73][29] = -8'd29;
        rom[73][30] = 8'd20;
        rom[73][31] = 8'd3;
        rom[74][0] = -8'd7;
        rom[74][1] = 8'd13;
        rom[74][2] = -8'd32;
        rom[74][3] = 8'd47;
        rom[74][4] = -8'd32;
        rom[74][5] = -8'd96;
        rom[74][6] = -8'd34;
        rom[74][7] = 8'd28;
        rom[74][8] = 8'd11;
        rom[74][9] = 8'd7;
        rom[74][10] = 8'd15;
        rom[74][11] = 8'd20;
        rom[74][12] = 8'd34;
        rom[74][13] = 8'd4;
        rom[74][14] = 8'd40;
        rom[74][15] = 8'd20;
        rom[74][16] = 8'd18;
        rom[74][17] = -8'd25;
        rom[74][18] = 8'd15;
        rom[74][19] = 8'd69;
        rom[74][20] = -8'd33;
        rom[74][21] = -8'd64;
        rom[74][22] = 8'd20;
        rom[74][23] = 8'd27;
        rom[74][24] = -8'd80;
        rom[74][25] = 8'd1;
        rom[74][26] = 8'd13;
        rom[74][27] = 8'd72;
        rom[74][28] = 8'd9;
        rom[74][29] = -8'd6;
        rom[74][30] = -8'd11;
        rom[74][31] = 8'd3;
        rom[75][0] = -8'd42;
        rom[75][1] = -8'd5;
        rom[75][2] = -8'd49;
        rom[75][3] = -8'd28;
        rom[75][4] = -8'd18;
        rom[75][5] = 8'd5;
        rom[75][6] = 8'd20;
        rom[75][7] = 8'd39;
        rom[75][8] = -8'd18;
        rom[75][9] = -8'd4;
        rom[75][10] = 8'd3;
        rom[75][11] = 8'd14;
        rom[75][12] = -8'd25;
        rom[75][13] = -8'd22;
        rom[75][14] = -8'd9;
        rom[75][15] = 8'd3;
        rom[75][16] = 8'd17;
        rom[75][17] = -8'd22;
        rom[75][18] = -8'd44;
        rom[75][19] = -8'd38;
        rom[75][20] = -8'd5;
        rom[75][21] = 8'd31;
        rom[75][22] = 8'd5;
        rom[75][23] = -8'd13;
        rom[75][24] = 8'd13;
        rom[75][25] = 8'd29;
        rom[75][26] = -8'd4;
        rom[75][27] = 8'd21;
        rom[75][28] = -8'd44;
        rom[75][29] = 8'd15;
        rom[75][30] = 8'd29;
        rom[75][31] = -8'd14;
        rom[76][0] = 8'd36;
        rom[76][1] = 8'd1;
        rom[76][2] = 8'd12;
        rom[76][3] = 8'd4;
        rom[76][4] = -8'd16;
        rom[76][5] = -8'd2;
        rom[76][6] = 8'd7;
        rom[76][7] = 8'd33;
        rom[76][8] = 8'd15;
        rom[76][9] = 8'd32;
        rom[76][10] = 8'd1;
        rom[76][11] = 8'd10;
        rom[76][12] = -8'd55;
        rom[76][13] = -8'd10;
        rom[76][14] = -8'd5;
        rom[76][15] = 8'd14;
        rom[76][16] = 8'd46;
        rom[76][17] = -8'd2;
        rom[76][18] = -8'd14;
        rom[76][19] = -8'd45;
        rom[76][20] = 8'd19;
        rom[76][21] = 8'd8;
        rom[76][22] = -8'd13;
        rom[76][23] = -8'd18;
        rom[76][24] = -8'd7;
        rom[76][25] = -8'd16;
        rom[76][26] = -8'd15;
        rom[76][27] = 8'd24;
        rom[76][28] = -8'd31;
        rom[76][29] = 8'd9;
        rom[76][30] = 8'd58;
        rom[76][31] = -8'd13;
        rom[77][0] = -8'd6;
        rom[77][1] = 8'd18;
        rom[77][2] = -8'd20;
        rom[77][3] = -8'd56;
        rom[77][4] = 8'd42;
        rom[77][5] = -8'd36;
        rom[77][6] = 8'd34;
        rom[77][7] = 8'd13;
        rom[77][8] = -8'd32;
        rom[77][9] = 8'd14;
        rom[77][10] = -8'd52;
        rom[77][11] = -8'd11;
        rom[77][12] = -8'd24;
        rom[77][13] = -8'd5;
        rom[77][14] = 8'd19;
        rom[77][15] = 8'd16;
        rom[77][16] = 8'd13;
        rom[77][17] = 8'd21;
        rom[77][18] = 8'd9;
        rom[77][19] = 8'd22;
        rom[77][20] = -8'd23;
        rom[77][21] = 8'd5;
        rom[77][22] = 8'd27;
        rom[77][23] = 8'd46;
        rom[77][24] = -8'd2;
        rom[77][25] = 8'd7;
        rom[77][26] = -8'd15;
        rom[77][27] = -8'd3;
        rom[77][28] = -8'd40;
        rom[77][29] = 8'd12;
        rom[77][30] = -8'd28;
        rom[77][31] = -8'd19;
        rom[78][0] = -8'd34;
        rom[78][1] = 8'd30;
        rom[78][2] = -8'd15;
        rom[78][3] = 8'd21;
        rom[78][4] = 8'd28;
        rom[78][5] = 8'd41;
        rom[78][6] = 8'd14;
        rom[78][7] = 8'd3;
        rom[78][8] = 8'd5;
        rom[78][9] = -8'd13;
        rom[78][10] = -8'd34;
        rom[78][11] = 8'd17;
        rom[78][12] = 8'd49;
        rom[78][13] = 8'd36;
        rom[78][14] = -8'd10;
        rom[78][15] = -8'd20;
        rom[78][16] = -8'd4;
        rom[78][17] = 8'd8;
        rom[78][18] = -8'd19;
        rom[78][19] = 8'd12;
        rom[78][20] = -8'd19;
        rom[78][21] = 8'd61;
        rom[78][22] = -8'd1;
        rom[78][23] = -8'd20;
        rom[78][24] = 8'd14;
        rom[78][25] = 8'd26;
        rom[78][26] = 8'd31;
        rom[78][27] = -8'd37;
        rom[78][28] = -8'd5;
        rom[78][29] = 8'd4;
        rom[78][30] = 8'd20;
        rom[78][31] = -8'd10;
        rom[79][0] = -8'd43;
        rom[79][1] = 8'd11;
        rom[79][2] = -8'd128;
        rom[79][3] = 8'd1;
        rom[79][4] = 8'd46;
        rom[79][5] = -8'd32;
        rom[79][6] = -8'd2;
        rom[79][7] = 8'd50;
        rom[79][8] = -8'd4;
        rom[79][9] = -8'd1;
        rom[79][10] = -8'd23;
        rom[79][11] = 8'd6;
        rom[79][12] = -8'd11;
        rom[79][13] = -8'd80;
        rom[79][14] = 8'd35;
        rom[79][15] = -8'd33;
        rom[79][16] = 8'd21;
        rom[79][17] = -8'd31;
        rom[79][18] = -8'd89;
        rom[79][19] = 8'd34;
        rom[79][20] = 8'd9;
        rom[79][21] = 8'd39;
        rom[79][22] = 8'd24;
        rom[79][23] = 8'd15;
        rom[79][24] = 8'd17;
        rom[79][25] = -8'd15;
        rom[79][26] = -8'd11;
        rom[79][27] = 8'd56;
        rom[79][28] = -8'd27;
        rom[79][29] = -8'd1;
        rom[79][30] = 8'd9;
        rom[79][31] = 8'd10;
        rom[80][0] = -8'd31;
        rom[80][1] = -8'd60;
        rom[80][2] = 8'd25;
        rom[80][3] = -8'd111;
        rom[80][4] = -8'd16;
        rom[80][5] = 8'd5;
        rom[80][6] = -8'd3;
        rom[80][7] = 8'd2;
        rom[80][8] = -8'd31;
        rom[80][9] = -8'd2;
        rom[80][10] = -8'd3;
        rom[80][11] = 8'd5;
        rom[80][12] = -8'd16;
        rom[80][13] = -8'd11;
        rom[80][14] = -8'd2;
        rom[80][15] = -8'd14;
        rom[80][16] = -8'd3;
        rom[80][17] = 8'd33;
        rom[80][18] = -8'd35;
        rom[80][19] = 8'd17;
        rom[80][20] = 8'd6;
        rom[80][21] = 8'd11;
        rom[80][22] = -8'd8;
        rom[80][23] = 8'd16;
        rom[80][24] = -8'd50;
        rom[80][25] = -8'd5;
        rom[80][26] = -8'd21;
        rom[80][27] = -8'd36;
        rom[80][28] = 8'd22;
        rom[80][29] = 8'd49;
        rom[80][30] = -8'd46;
        rom[80][31] = 8'd7;
        rom[81][0] = 8'd1;
        rom[81][1] = -8'd2;
        rom[81][2] = -8'd22;
        rom[81][3] = 8'd39;
        rom[81][4] = -8'd51;
        rom[81][5] = 8'd8;
        rom[81][6] = 8'd12;
        rom[81][7] = -8'd2;
        rom[81][8] = 8'd23;
        rom[81][9] = -8'd2;
        rom[81][10] = 8'd29;
        rom[81][11] = 8'd13;
        rom[81][12] = 8'd5;
        rom[81][13] = -8'd21;
        rom[81][14] = -8'd7;
        rom[81][15] = -8'd3;
        rom[81][16] = 8'd3;
        rom[81][17] = -8'd30;
        rom[81][18] = 8'd12;
        rom[81][19] = 8'd17;
        rom[81][20] = 8'd27;
        rom[81][21] = -8'd15;
        rom[81][22] = -8'd54;
        rom[81][23] = -8'd8;
        rom[81][24] = 8'd20;
        rom[81][25] = 8'd11;
        rom[81][26] = 8'd18;
        rom[81][27] = 8'd35;
        rom[81][28] = -8'd17;
        rom[81][29] = -8'd6;
        rom[81][30] = 8'd11;
        rom[81][31] = -8'd13;
        rom[82][0] = -8'd22;
        rom[82][1] = -8'd10;
        rom[82][2] = -8'd12;
        rom[82][3] = 8'd22;
        rom[82][4] = -8'd25;
        rom[82][5] = 8'd7;
        rom[82][6] = -8'd53;
        rom[82][7] = 8'd22;
        rom[82][8] = 8'd20;
        rom[82][9] = -8'd35;
        rom[82][10] = -8'd1;
        rom[82][11] = 8'd13;
        rom[82][12] = -8'd59;
        rom[82][13] = 8'd4;
        rom[82][14] = 8'd10;
        rom[82][15] = -8'd50;
        rom[82][16] = 8'd20;
        rom[82][17] = -8'd26;
        rom[82][18] = 8'd13;
        rom[82][19] = 8'd36;
        rom[82][20] = 8'd5;
        rom[82][21] = -8'd29;
        rom[82][22] = 8'd23;
        rom[82][23] = -8'd33;
        rom[82][24] = -8'd8;
        rom[82][25] = 8'd19;
        rom[82][26] = -8'd10;
        rom[82][27] = -8'd5;
        rom[82][28] = -8'd1;
        rom[82][29] = 8'd6;
        rom[82][30] = 8'd26;
        rom[82][31] = 8'd28;
        rom[83][0] = -8'd1;
        rom[83][1] = -8'd61;
        rom[83][2] = 8'd2;
        rom[83][3] = -8'd10;
        rom[83][4] = -8'd51;
        rom[83][5] = 8'd5;
        rom[83][6] = 8'd33;
        rom[83][7] = -8'd14;
        rom[83][8] = -8'd23;
        rom[83][9] = 8'd13;
        rom[83][10] = 8'd35;
        rom[83][11] = 8'd38;
        rom[83][12] = 8'd62;
        rom[83][13] = -8'd24;
        rom[83][14] = -8'd48;
        rom[83][15] = -8'd35;
        rom[83][16] = 8'd19;
        rom[83][17] = -8'd8;
        rom[83][18] = -8'd11;
        rom[83][19] = -8'd2;
        rom[83][20] = 8'd19;
        rom[83][21] = -8'd1;
        rom[83][22] = 8'd35;
        rom[83][23] = -8'd30;
        rom[83][24] = -8'd16;
        rom[83][25] = 8'd6;
        rom[83][26] = -8'd38;
        rom[83][27] = -8'd28;
        rom[83][28] = 8'd30;
        rom[83][29] = -8'd21;
        rom[83][30] = 8'd25;
        rom[83][31] = 8'd8;
        rom[84][0] = -8'd3;
        rom[84][1] = -8'd25;
        rom[84][2] = 8'd11;
        rom[84][3] = -8'd33;
        rom[84][4] = -8'd23;
        rom[84][5] = 8'd5;
        rom[84][6] = 8'd7;
        rom[84][7] = -8'd16;
        rom[84][8] = -8'd23;
        rom[84][9] = 8'd21;
        rom[84][10] = 8'd10;
        rom[84][11] = 8'd59;
        rom[84][12] = -8'd5;
        rom[84][13] = 8'd34;
        rom[84][14] = 8'd12;
        rom[84][15] = -8'd27;
        rom[84][16] = 8'd7;
        rom[84][17] = 8'd37;
        rom[84][18] = -8'd8;
        rom[84][19] = 8'd1;
        rom[84][20] = 8'd17;
        rom[84][21] = 8'd27;
        rom[84][22] = 8'd20;
        rom[84][23] = -8'd7;
        rom[84][24] = -8'd3;
        rom[84][25] = -8'd7;
        rom[84][26] = -8'd9;
        rom[84][27] = 8'd18;
        rom[84][28] = 8'd10;
        rom[84][29] = -8'd36;
        rom[84][30] = 8'd16;
        rom[84][31] = 8'd22;
        rom[85][0] = 8'd9;
        rom[85][1] = -8'd21;
        rom[85][2] = -8'd67;
        rom[85][3] = -8'd2;
        rom[85][4] = -8'd66;
        rom[85][5] = 8'd3;
        rom[85][6] = 8'd19;
        rom[85][7] = 8'd22;
        rom[85][8] = -8'd7;
        rom[85][9] = -8'd85;
        rom[85][10] = 8'd33;
        rom[85][11] = 8'd18;
        rom[85][12] = -8'd57;
        rom[85][13] = -8'd33;
        rom[85][14] = -8'd3;
        rom[85][15] = 8'd19;
        rom[85][16] = -8'd8;
        rom[85][17] = 8'd19;
        rom[85][18] = -8'd48;
        rom[85][19] = -8'd42;
        rom[85][20] = -8'd11;
        rom[85][21] = 8'd3;
        rom[85][22] = 8'd39;
        rom[85][23] = 8'd22;
        rom[85][24] = -8'd10;
        rom[85][25] = 8'd49;
        rom[85][26] = -8'd6;
        rom[85][27] = -8'd5;
        rom[85][28] = 8'd36;
        rom[85][29] = 8'd7;
        rom[85][30] = -8'd9;
        rom[85][31] = 8'd15;
        rom[86][0] = 8'd13;
        rom[86][1] = -8'd39;
        rom[86][2] = 8'd7;
        rom[86][3] = -8'd13;
        rom[86][4] = 8'd31;
        rom[86][5] = -8'd47;
        rom[86][6] = -8'd8;
        rom[86][7] = -8'd13;
        rom[86][8] = -8'd6;
        rom[86][9] = 8'd24;
        rom[86][10] = -8'd34;
        rom[86][11] = 8'd18;
        rom[86][12] = -8'd4;
        rom[86][13] = 8'd7;
        rom[86][14] = 8'd29;
        rom[86][15] = -8'd29;
        rom[86][16] = -8'd22;
        rom[86][17] = -8'd5;
        rom[86][18] = 8'd20;
        rom[86][19] = 8'd29;
        rom[86][20] = 8'd2;
        rom[86][21] = -8'd4;
        rom[86][22] = -8'd15;
        rom[86][23] = -8'd2;
        rom[86][24] = 8'd19;
        rom[86][25] = -8'd54;
        rom[86][26] = -8'd8;
        rom[86][27] = -8'd6;
        rom[86][28] = 8'd19;
        rom[86][29] = 8'd46;
        rom[86][30] = 8'd19;
        rom[86][31] = 8'd27;
        rom[87][0] = 8'd24;
        rom[87][1] = -8'd47;
        rom[87][2] = -8'd37;
        rom[87][3] = -8'd31;
        rom[87][4] = -8'd41;
        rom[87][5] = -8'd31;
        rom[87][6] = 8'd37;
        rom[87][7] = 8'd39;
        rom[87][8] = 8'd2;
        rom[87][9] = -8'd10;
        rom[87][10] = 8'd63;
        rom[87][11] = 8'd2;
        rom[87][12] = -8'd48;
        rom[87][13] = -8'd52;
        rom[87][14] = -8'd1;
        rom[87][15] = 8'd18;
        rom[87][16] = 8'd22;
        rom[87][17] = 8'd23;
        rom[87][18] = -8'd20;
        rom[87][19] = 8'd0;
        rom[87][20] = 8'd3;
        rom[87][21] = -8'd31;
        rom[87][22] = 8'd24;
        rom[87][23] = 8'd13;
        rom[87][24] = 8'd0;
        rom[87][25] = 8'd13;
        rom[87][26] = -8'd14;
        rom[87][27] = 8'd16;
        rom[87][28] = 8'd12;
        rom[87][29] = 8'd16;
        rom[87][30] = 8'd4;
        rom[87][31] = 8'd28;
        rom[88][0] = 8'd11;
        rom[88][1] = -8'd23;
        rom[88][2] = 8'd21;
        rom[88][3] = -8'd18;
        rom[88][4] = -8'd13;
        rom[88][5] = -8'd18;
        rom[88][6] = 8'd12;
        rom[88][7] = 8'd1;
        rom[88][8] = -8'd1;
        rom[88][9] = -8'd2;
        rom[88][10] = -8'd10;
        rom[88][11] = 8'd38;
        rom[88][12] = -8'd16;
        rom[88][13] = 8'd26;
        rom[88][14] = 8'd24;
        rom[88][15] = 8'd33;
        rom[88][16] = -8'd51;
        rom[88][17] = 8'd45;
        rom[88][18] = 8'd4;
        rom[88][19] = -8'd67;
        rom[88][20] = -8'd64;
        rom[88][21] = 8'd7;
        rom[88][22] = 8'd19;
        rom[88][23] = 8'd21;
        rom[88][24] = -8'd51;
        rom[88][25] = -8'd16;
        rom[88][26] = 8'd8;
        rom[88][27] = 8'd1;
        rom[88][28] = 8'd32;
        rom[88][29] = -8'd10;
        rom[88][30] = -8'd24;
        rom[88][31] = 8'd20;
        rom[89][0] = -8'd5;
        rom[89][1] = -8'd4;
        rom[89][2] = 8'd14;
        rom[89][3] = 8'd20;
        rom[89][4] = 8'd23;
        rom[89][5] = 8'd12;
        rom[89][6] = -8'd9;
        rom[89][7] = -8'd27;
        rom[89][8] = -8'd36;
        rom[89][9] = -8'd6;
        rom[89][10] = 8'd18;
        rom[89][11] = 8'd21;
        rom[89][12] = 8'd22;
        rom[89][13] = -8'd38;
        rom[89][14] = -8'd12;
        rom[89][15] = 8'd32;
        rom[89][16] = -8'd1;
        rom[89][17] = 8'd22;
        rom[89][18] = 8'd1;
        rom[89][19] = 8'd0;
        rom[89][20] = -8'd38;
        rom[89][21] = -8'd19;
        rom[89][22] = 8'd3;
        rom[89][23] = 8'd11;
        rom[89][24] = -8'd33;
        rom[89][25] = 8'd14;
        rom[89][26] = 8'd25;
        rom[89][27] = -8'd23;
        rom[89][28] = -8'd7;
        rom[89][29] = 8'd2;
        rom[89][30] = -8'd33;
        rom[89][31] = 8'd19;
        rom[90][0] = 8'd6;
        rom[90][1] = -8'd20;
        rom[90][2] = -8'd47;
        rom[90][3] = 8'd33;
        rom[90][4] = -8'd17;
        rom[90][5] = -8'd90;
        rom[90][6] = -8'd47;
        rom[90][7] = 8'd25;
        rom[90][8] = 8'd14;
        rom[90][9] = 8'd15;
        rom[90][10] = 8'd18;
        rom[90][11] = 8'd19;
        rom[90][12] = -8'd9;
        rom[90][13] = 8'd31;
        rom[90][14] = 8'd21;
        rom[90][15] = -8'd22;
        rom[90][16] = 8'd20;
        rom[90][17] = -8'd7;
        rom[90][18] = 8'd26;
        rom[90][19] = 8'd40;
        rom[90][20] = -8'd12;
        rom[90][21] = -8'd43;
        rom[90][22] = 8'd49;
        rom[90][23] = 8'd5;
        rom[90][24] = -8'd5;
        rom[90][25] = -8'd46;
        rom[90][26] = 8'd18;
        rom[90][27] = 8'd38;
        rom[90][28] = -8'd1;
        rom[90][29] = 8'd0;
        rom[90][30] = 8'd45;
        rom[90][31] = 8'd23;
        rom[91][0] = 8'd14;
        rom[91][1] = 8'd6;
        rom[91][2] = -8'd50;
        rom[91][3] = 8'd11;
        rom[91][4] = -8'd40;
        rom[91][5] = -8'd20;
        rom[91][6] = -8'd16;
        rom[91][7] = 8'd1;
        rom[91][8] = -8'd15;
        rom[91][9] = -8'd21;
        rom[91][10] = 8'd17;
        rom[91][11] = -8'd9;
        rom[91][12] = -8'd7;
        rom[91][13] = -8'd19;
        rom[91][14] = -8'd8;
        rom[91][15] = 8'd26;
        rom[91][16] = 8'd2;
        rom[91][17] = -8'd17;
        rom[91][18] = -8'd48;
        rom[91][19] = -8'd19;
        rom[91][20] = -8'd9;
        rom[91][21] = 8'd18;
        rom[91][22] = 8'd7;
        rom[91][23] = -8'd33;
        rom[91][24] = -8'd8;
        rom[91][25] = 8'd21;
        rom[91][26] = 8'd4;
        rom[91][27] = -8'd11;
        rom[91][28] = 8'd20;
        rom[91][29] = -8'd21;
        rom[91][30] = -8'd2;
        rom[91][31] = 8'd15;
        rom[92][0] = 8'd41;
        rom[92][1] = 8'd2;
        rom[92][2] = 8'd24;
        rom[92][3] = -8'd5;
        rom[92][4] = 8'd33;
        rom[92][5] = -8'd51;
        rom[92][6] = 8'd29;
        rom[92][7] = 8'd24;
        rom[92][8] = 8'd25;
        rom[92][9] = 8'd15;
        rom[92][10] = 8'd18;
        rom[92][11] = 8'd8;
        rom[92][12] = -8'd66;
        rom[92][13] = -8'd15;
        rom[92][14] = 8'd4;
        rom[92][15] = -8'd19;
        rom[92][16] = 8'd17;
        rom[92][17] = -8'd4;
        rom[92][18] = -8'd1;
        rom[92][19] = -8'd29;
        rom[92][20] = -8'd30;
        rom[92][21] = 8'd2;
        rom[92][22] = -8'd25;
        rom[92][23] = -8'd13;
        rom[92][24] = -8'd9;
        rom[92][25] = 8'd37;
        rom[92][26] = -8'd5;
        rom[92][27] = -8'd14;
        rom[92][28] = -8'd31;
        rom[92][29] = -8'd3;
        rom[92][30] = -8'd15;
        rom[92][31] = -8'd10;
        rom[93][0] = 8'd5;
        rom[93][1] = 8'd6;
        rom[93][2] = -8'd11;
        rom[93][3] = -8'd29;
        rom[93][4] = 8'd47;
        rom[93][5] = -8'd16;
        rom[93][6] = 8'd3;
        rom[93][7] = -8'd14;
        rom[93][8] = -8'd7;
        rom[93][9] = -8'd22;
        rom[93][10] = 8'd11;
        rom[93][11] = -8'd11;
        rom[93][12] = -8'd50;
        rom[93][13] = -8'd11;
        rom[93][14] = -8'd18;
        rom[93][15] = -8'd5;
        rom[93][16] = 8'd5;
        rom[93][17] = 8'd17;
        rom[93][18] = 8'd14;
        rom[93][19] = 8'd6;
        rom[93][20] = -8'd8;
        rom[93][21] = -8'd35;
        rom[93][22] = 8'd15;
        rom[93][23] = 8'd1;
        rom[93][24] = 8'd5;
        rom[93][25] = 8'd19;
        rom[93][26] = 8'd20;
        rom[93][27] = -8'd6;
        rom[93][28] = 8'd2;
        rom[93][29] = -8'd13;
        rom[93][30] = -8'd48;
        rom[93][31] = 8'd4;
        rom[94][0] = -8'd18;
        rom[94][1] = 8'd56;
        rom[94][2] = -8'd36;
        rom[94][3] = 8'd18;
        rom[94][4] = -8'd34;
        rom[94][5] = 8'd16;
        rom[94][6] = -8'd33;
        rom[94][7] = -8'd3;
        rom[94][8] = 8'd23;
        rom[94][9] = -8'd39;
        rom[94][10] = -8'd9;
        rom[94][11] = 8'd33;
        rom[94][12] = 8'd42;
        rom[94][13] = -8'd37;
        rom[94][14] = -8'd4;
        rom[94][15] = -8'd21;
        rom[94][16] = 8'd9;
        rom[94][17] = -8'd41;
        rom[94][18] = 8'd8;
        rom[94][19] = 8'd14;
        rom[94][20] = 8'd17;
        rom[94][21] = 8'd24;
        rom[94][22] = -8'd6;
        rom[94][23] = -8'd13;
        rom[94][24] = 8'd14;
        rom[94][25] = -8'd6;
        rom[94][26] = -8'd13;
        rom[94][27] = -8'd20;
        rom[94][28] = 8'd5;
        rom[94][29] = 8'd7;
        rom[94][30] = -8'd14;
        rom[94][31] = -8'd12;
        rom[95][0] = -8'd9;
        rom[95][1] = -8'd21;
        rom[95][2] = -8'd128;
        rom[95][3] = -8'd20;
        rom[95][4] = 8'd13;
        rom[95][5] = -8'd28;
        rom[95][6] = -8'd8;
        rom[95][7] = 8'd28;
        rom[95][8] = 8'd22;
        rom[95][9] = -8'd22;
        rom[95][10] = -8'd15;
        rom[95][11] = 8'd4;
        rom[95][12] = 8'd5;
        rom[95][13] = -8'd50;
        rom[95][14] = -8'd3;
        rom[95][15] = -8'd33;
        rom[95][16] = 8'd29;
        rom[95][17] = -8'd12;
        rom[95][18] = -8'd7;
        rom[95][19] = 8'd25;
        rom[95][20] = 8'd9;
        rom[95][21] = -8'd9;
        rom[95][22] = 8'd14;
        rom[95][23] = -8'd22;
        rom[95][24] = 8'd25;
        rom[95][25] = 8'd12;
        rom[95][26] = 8'd4;
        rom[95][27] = -8'd15;
        rom[95][28] = 8'd2;
        rom[95][29] = 8'd15;
        rom[95][30] = 8'd27;
        rom[95][31] = 8'd14;
        rom[96][0] = -8'd9;
        rom[96][1] = 8'd38;
        rom[96][2] = 8'd26;
        rom[96][3] = -8'd33;
        rom[96][4] = -8'd18;
        rom[96][5] = 8'd8;
        rom[96][6] = -8'd18;
        rom[96][7] = 8'd19;
        rom[96][8] = 8'd30;
        rom[96][9] = 8'd15;
        rom[96][10] = 8'd6;
        rom[96][11] = -8'd22;
        rom[96][12] = -8'd12;
        rom[96][13] = 8'd9;
        rom[96][14] = -8'd3;
        rom[96][15] = -8'd20;
        rom[96][16] = -8'd21;
        rom[96][17] = 8'd4;
        rom[96][18] = 8'd12;
        rom[96][19] = 8'd35;
        rom[96][20] = 8'd12;
        rom[96][21] = 8'd9;
        rom[96][22] = 8'd0;
        rom[96][23] = -8'd27;
        rom[96][24] = 8'd32;
        rom[96][25] = 8'd21;
        rom[96][26] = -8'd18;
        rom[96][27] = 8'd10;
        rom[96][28] = 8'd12;
        rom[96][29] = 8'd12;
        rom[96][30] = -8'd53;
        rom[96][31] = 8'd3;
        rom[97][0] = -8'd17;
        rom[97][1] = -8'd4;
        rom[97][2] = -8'd8;
        rom[97][3] = -8'd25;
        rom[97][4] = 8'd9;
        rom[97][5] = -8'd2;
        rom[97][6] = -8'd24;
        rom[97][7] = -8'd12;
        rom[97][8] = -8'd17;
        rom[97][9] = 8'd16;
        rom[97][10] = -8'd23;
        rom[97][11] = 8'd0;
        rom[97][12] = -8'd18;
        rom[97][13] = 8'd37;
        rom[97][14] = -8'd34;
        rom[97][15] = -8'd26;
        rom[97][16] = 8'd12;
        rom[97][17] = 8'd9;
        rom[97][18] = -8'd19;
        rom[97][19] = 8'd21;
        rom[97][20] = -8'd38;
        rom[97][21] = -8'd11;
        rom[97][22] = -8'd3;
        rom[97][23] = 8'd10;
        rom[97][24] = 8'd19;
        rom[97][25] = -8'd16;
        rom[97][26] = -8'd30;
        rom[97][27] = 8'd25;
        rom[97][28] = -8'd10;
        rom[97][29] = 8'd1;
        rom[97][30] = -8'd5;
        rom[97][31] = 8'd22;
        rom[98][0] = 8'd11;
        rom[98][1] = 8'd45;
        rom[98][2] = 8'd19;
        rom[98][3] = -8'd15;
        rom[98][4] = -8'd28;
        rom[98][5] = -8'd9;
        rom[98][6] = 8'd37;
        rom[98][7] = 8'd13;
        rom[98][8] = -8'd14;
        rom[98][9] = 8'd0;
        rom[98][10] = -8'd50;
        rom[98][11] = -8'd11;
        rom[98][12] = 8'd42;
        rom[98][13] = 8'd22;
        rom[98][14] = 8'd21;
        rom[98][15] = -8'd13;
        rom[98][16] = 8'd5;
        rom[98][17] = 8'd11;
        rom[98][18] = -8'd19;
        rom[98][19] = -8'd6;
        rom[98][20] = -8'd13;
        rom[98][21] = 8'd15;
        rom[98][22] = -8'd51;
        rom[98][23] = 8'd8;
        rom[98][24] = -8'd1;
        rom[98][25] = 8'd22;
        rom[98][26] = 8'd5;
        rom[98][27] = -8'd4;
        rom[98][28] = -8'd13;
        rom[98][29] = -8'd37;
        rom[98][30] = 8'd8;
        rom[98][31] = -8'd42;
        rom[99][0] = 8'd9;
        rom[99][1] = 8'd64;
        rom[99][2] = 8'd14;
        rom[99][3] = -8'd20;
        rom[99][4] = 8'd16;
        rom[99][5] = -8'd12;
        rom[99][6] = -8'd32;
        rom[99][7] = 8'd15;
        rom[99][8] = 8'd35;
        rom[99][9] = -8'd9;
        rom[99][10] = -8'd21;
        rom[99][11] = -8'd27;
        rom[99][12] = -8'd33;
        rom[99][13] = -8'd4;
        rom[99][14] = 8'd31;
        rom[99][15] = 8'd14;
        rom[99][16] = -8'd4;
        rom[99][17] = 8'd0;
        rom[99][18] = -8'd22;
        rom[99][19] = 8'd10;
        rom[99][20] = 8'd11;
        rom[99][21] = 8'd1;
        rom[99][22] = 8'd9;
        rom[99][23] = 8'd23;
        rom[99][24] = 8'd6;
        rom[99][25] = -8'd8;
        rom[99][26] = -8'd45;
        rom[99][27] = 8'd22;
        rom[99][28] = -8'd35;
        rom[99][29] = 8'd15;
        rom[99][30] = -8'd52;
        rom[99][31] = 8'd8;
        rom[100][0] = 8'd37;
        rom[100][1] = 8'd23;
        rom[100][2] = -8'd9;
        rom[100][3] = -8'd11;
        rom[100][4] = -8'd4;
        rom[100][5] = -8'd31;
        rom[100][6] = -8'd27;
        rom[100][7] = -8'd11;
        rom[100][8] = 8'd22;
        rom[100][9] = 8'd2;
        rom[100][10] = -8'd6;
        rom[100][11] = -8'd49;
        rom[100][12] = -8'd1;
        rom[100][13] = 8'd2;
        rom[100][14] = 8'd10;
        rom[100][15] = -8'd17;
        rom[100][16] = -8'd55;
        rom[100][17] = 8'd24;
        rom[100][18] = -8'd1;
        rom[100][19] = 8'd21;
        rom[100][20] = -8'd70;
        rom[100][21] = 8'd10;
        rom[100][22] = -8'd7;
        rom[100][23] = -8'd17;
        rom[100][24] = 8'd17;
        rom[100][25] = 8'd11;
        rom[100][26] = 8'd12;
        rom[100][27] = 8'd0;
        rom[100][28] = -8'd32;
        rom[100][29] = -8'd15;
        rom[100][30] = -8'd21;
        rom[100][31] = -8'd8;
        rom[101][0] = 8'd23;
        rom[101][1] = 8'd17;
        rom[101][2] = 8'd3;
        rom[101][3] = 8'd33;
        rom[101][4] = 8'd6;
        rom[101][5] = -8'd2;
        rom[101][6] = -8'd19;
        rom[101][7] = 8'd16;
        rom[101][8] = -8'd5;
        rom[101][9] = 8'd0;
        rom[101][10] = -8'd19;
        rom[101][11] = 8'd4;
        rom[101][12] = 8'd20;
        rom[101][13] = 8'd17;
        rom[101][14] = 8'd26;
        rom[101][15] = -8'd3;
        rom[101][16] = 8'd24;
        rom[101][17] = 8'd0;
        rom[101][18] = -8'd8;
        rom[101][19] = -8'd13;
        rom[101][20] = 8'd5;
        rom[101][21] = 8'd9;
        rom[101][22] = 8'd26;
        rom[101][23] = -8'd14;
        rom[101][24] = -8'd19;
        rom[101][25] = 8'd9;
        rom[101][26] = 8'd3;
        rom[101][27] = -8'd29;
        rom[101][28] = 8'd4;
        rom[101][29] = 8'd17;
        rom[101][30] = -8'd15;
        rom[101][31] = -8'd128;
        rom[102][0] = 8'd1;
        rom[102][1] = -8'd12;
        rom[102][2] = -8'd21;
        rom[102][3] = 8'd1;
        rom[102][4] = -8'd13;
        rom[102][5] = 8'd0;
        rom[102][6] = -8'd3;
        rom[102][7] = 8'd15;
        rom[102][8] = 8'd32;
        rom[102][9] = -8'd2;
        rom[102][10] = 8'd7;
        rom[102][11] = -8'd22;
        rom[102][12] = -8'd4;
        rom[102][13] = 8'd10;
        rom[102][14] = -8'd19;
        rom[102][15] = 8'd14;
        rom[102][16] = -8'd14;
        rom[102][17] = -8'd6;
        rom[102][18] = 8'd31;
        rom[102][19] = -8'd4;
        rom[102][20] = 8'd17;
        rom[102][21] = 8'd11;
        rom[102][22] = -8'd32;
        rom[102][23] = 8'd20;
        rom[102][24] = 8'd26;
        rom[102][25] = -8'd8;
        rom[102][26] = 8'd11;
        rom[102][27] = 8'd3;
        rom[102][28] = -8'd15;
        rom[102][29] = 8'd10;
        rom[102][30] = 8'd36;
        rom[102][31] = 8'd7;
        rom[103][0] = 8'd28;
        rom[103][1] = 8'd23;
        rom[103][2] = 8'd35;
        rom[103][3] = 8'd5;
        rom[103][4] = 8'd33;
        rom[103][5] = 8'd9;
        rom[103][6] = 8'd3;
        rom[103][7] = -8'd4;
        rom[103][8] = -8'd33;
        rom[103][9] = -8'd18;
        rom[103][10] = 8'd4;
        rom[103][11] = -8'd1;
        rom[103][12] = 8'd17;
        rom[103][13] = -8'd5;
        rom[103][14] = -8'd14;
        rom[103][15] = -8'd15;
        rom[103][16] = -8'd10;
        rom[103][17] = 8'd18;
        rom[103][18] = 8'd1;
        rom[103][19] = 8'd28;
        rom[103][20] = 8'd14;
        rom[103][21] = -8'd31;
        rom[103][22] = 8'd27;
        rom[103][23] = 8'd17;
        rom[103][24] = 8'd20;
        rom[103][25] = -8'd15;
        rom[103][26] = 8'd0;
        rom[103][27] = -8'd10;
        rom[103][28] = -8'd5;
        rom[103][29] = -8'd14;
        rom[103][30] = 8'd1;
        rom[103][31] = -8'd22;
        rom[104][0] = 8'd6;
        rom[104][1] = 8'd14;
        rom[104][2] = 8'd21;
        rom[104][3] = -8'd33;
        rom[104][4] = -8'd8;
        rom[104][5] = -8'd33;
        rom[104][6] = 8'd26;
        rom[104][7] = -8'd3;
        rom[104][8] = 8'd11;
        rom[104][9] = 8'd23;
        rom[104][10] = 8'd2;
        rom[104][11] = -8'd48;
        rom[104][12] = 8'd14;
        rom[104][13] = -8'd18;
        rom[104][14] = -8'd17;
        rom[104][15] = 8'd19;
        rom[104][16] = -8'd67;
        rom[104][17] = 8'd16;
        rom[104][18] = 8'd13;
        rom[104][19] = -8'd27;
        rom[104][20] = -8'd45;
        rom[104][21] = 8'd9;
        rom[104][22] = -8'd5;
        rom[104][23] = 8'd26;
        rom[104][24] = -8'd2;
        rom[104][25] = 8'd6;
        rom[104][26] = 8'd41;
        rom[104][27] = 8'd6;
        rom[104][28] = 8'd19;
        rom[104][29] = 8'd4;
        rom[104][30] = 8'd15;
        rom[104][31] = 8'd3;
        rom[105][0] = -8'd7;
        rom[105][1] = -8'd13;
        rom[105][2] = 8'd12;
        rom[105][3] = -8'd27;
        rom[105][4] = -8'd6;
        rom[105][5] = -8'd10;
        rom[105][6] = 8'd0;
        rom[105][7] = 8'd15;
        rom[105][8] = -8'd51;
        rom[105][9] = 8'd40;
        rom[105][10] = 8'd1;
        rom[105][11] = -8'd13;
        rom[105][12] = -8'd35;
        rom[105][13] = 8'd1;
        rom[105][14] = 8'd6;
        rom[105][15] = -8'd7;
        rom[105][16] = -8'd19;
        rom[105][17] = 8'd11;
        rom[105][18] = 8'd33;
        rom[105][19] = 8'd5;
        rom[105][20] = -8'd29;
        rom[105][21] = -8'd9;
        rom[105][22] = 8'd15;
        rom[105][23] = -8'd3;
        rom[105][24] = -8'd2;
        rom[105][25] = -8'd3;
        rom[105][26] = 8'd5;
        rom[105][27] = 8'd19;
        rom[105][28] = -8'd5;
        rom[105][29] = -8'd7;
        rom[105][30] = 8'd13;
        rom[105][31] = 8'd13;
        rom[106][0] = 8'd3;
        rom[106][1] = 8'd32;
        rom[106][2] = 8'd10;
        rom[106][3] = -8'd4;
        rom[106][4] = -8'd12;
        rom[106][5] = 8'd4;
        rom[106][6] = -8'd2;
        rom[106][7] = -8'd9;
        rom[106][8] = -8'd22;
        rom[106][9] = 8'd37;
        rom[106][10] = 8'd11;
        rom[106][11] = 8'd19;
        rom[106][12] = 8'd15;
        rom[106][13] = 8'd26;
        rom[106][14] = -8'd24;
        rom[106][15] = -8'd30;
        rom[106][16] = -8'd3;
        rom[106][17] = 8'd13;
        rom[106][18] = 8'd14;
        rom[106][19] = -8'd4;
        rom[106][20] = -8'd33;
        rom[106][21] = 8'd4;
        rom[106][22] = 8'd5;
        rom[106][23] = 8'd13;
        rom[106][24] = 8'd20;
        rom[106][25] = 8'd27;
        rom[106][26] = -8'd1;
        rom[106][27] = -8'd9;
        rom[106][28] = 8'd28;
        rom[106][29] = -8'd25;
        rom[106][30] = -8'd16;
        rom[106][31] = 8'd3;
        rom[107][0] = 8'd28;
        rom[107][1] = 8'd28;
        rom[107][2] = -8'd4;
        rom[107][3] = 8'd38;
        rom[107][4] = 8'd9;
        rom[107][5] = 8'd16;
        rom[107][6] = -8'd10;
        rom[107][7] = 8'd22;
        rom[107][8] = 8'd20;
        rom[107][9] = -8'd7;
        rom[107][10] = -8'd47;
        rom[107][11] = 8'd21;
        rom[107][12] = 8'd12;
        rom[107][13] = 8'd56;
        rom[107][14] = 8'd14;
        rom[107][15] = -8'd15;
        rom[107][16] = -8'd41;
        rom[107][17] = 8'd1;
        rom[107][18] = -8'd54;
        rom[107][19] = -8'd6;
        rom[107][20] = 8'd34;
        rom[107][21] = 8'd28;
        rom[107][22] = -8'd3;
        rom[107][23] = -8'd11;
        rom[107][24] = 8'd24;
        rom[107][25] = -8'd10;
        rom[107][26] = 8'd22;
        rom[107][27] = -8'd8;
        rom[107][28] = 8'd10;
        rom[107][29] = -8'd7;
        rom[107][30] = 8'd30;
        rom[107][31] = -8'd56;
        rom[108][0] = 8'd13;
        rom[108][1] = 8'd0;
        rom[108][2] = 8'd2;
        rom[108][3] = -8'd20;
        rom[108][4] = -8'd22;
        rom[108][5] = -8'd2;
        rom[108][6] = 8'd2;
        rom[108][7] = 8'd7;
        rom[108][8] = 8'd14;
        rom[108][9] = -8'd15;
        rom[108][10] = -8'd32;
        rom[108][11] = -8'd33;
        rom[108][12] = 8'd26;
        rom[108][13] = -8'd7;
        rom[108][14] = 8'd3;
        rom[108][15] = 8'd25;
        rom[108][16] = 8'd4;
        rom[108][17] = 8'd3;
        rom[108][18] = 8'd27;
        rom[108][19] = -8'd1;
        rom[108][20] = 8'd12;
        rom[108][21] = -8'd31;
        rom[108][22] = 8'd19;
        rom[108][23] = -8'd32;
        rom[108][24] = 8'd11;
        rom[108][25] = -8'd68;
        rom[108][26] = 8'd13;
        rom[108][27] = -8'd4;
        rom[108][28] = -8'd19;
        rom[108][29] = 8'd10;
        rom[108][30] = 8'd37;
        rom[108][31] = -8'd8;
        rom[109][0] = 8'd2;
        rom[109][1] = 8'd5;
        rom[109][2] = 8'd5;
        rom[109][3] = 8'd22;
        rom[109][4] = -8'd50;
        rom[109][5] = 8'd33;
        rom[109][6] = 8'd15;
        rom[109][7] = 8'd14;
        rom[109][8] = 8'd9;
        rom[109][9] = 8'd22;
        rom[109][10] = -8'd17;
        rom[109][11] = -8'd12;
        rom[109][12] = 8'd24;
        rom[109][13] = -8'd14;
        rom[109][14] = 8'd4;
        rom[109][15] = -8'd8;
        rom[109][16] = -8'd2;
        rom[109][17] = 8'd7;
        rom[109][18] = 8'd0;
        rom[109][19] = -8'd9;
        rom[109][20] = 8'd35;
        rom[109][21] = 8'd28;
        rom[109][22] = -8'd12;
        rom[109][23] = -8'd7;
        rom[109][24] = -8'd11;
        rom[109][25] = -8'd15;
        rom[109][26] = -8'd22;
        rom[109][27] = 8'd6;
        rom[109][28] = -8'd10;
        rom[109][29] = 8'd1;
        rom[109][30] = 8'd15;
        rom[109][31] = -8'd23;
        rom[110][0] = 8'd13;
        rom[110][1] = -8'd16;
        rom[110][2] = -8'd8;
        rom[110][3] = -8'd30;
        rom[110][4] = -8'd36;
        rom[110][5] = -8'd3;
        rom[110][6] = -8'd24;
        rom[110][7] = -8'd6;
        rom[110][8] = 8'd3;
        rom[110][9] = 8'd27;
        rom[110][10] = -8'd6;
        rom[110][11] = 8'd6;
        rom[110][12] = -8'd30;
        rom[110][13] = 8'd13;
        rom[110][14] = 8'd29;
        rom[110][15] = -8'd17;
        rom[110][16] = -8'd12;
        rom[110][17] = -8'd4;
        rom[110][18] = -8'd21;
        rom[110][19] = 8'd4;
        rom[110][20] = -8'd8;
        rom[110][21] = 8'd5;
        rom[110][22] = 8'd2;
        rom[110][23] = -8'd31;
        rom[110][24] = -8'd11;
        rom[110][25] = -8'd4;
        rom[110][26] = 8'd13;
        rom[110][27] = 8'd22;
        rom[110][28] = 8'd24;
        rom[110][29] = 8'd27;
        rom[110][30] = 8'd10;
        rom[110][31] = -8'd24;
        rom[111][0] = 8'd1;
        rom[111][1] = 8'd10;
        rom[111][2] = -8'd34;
        rom[111][3] = 8'd17;
        rom[111][4] = -8'd20;
        rom[111][5] = 8'd23;
        rom[111][6] = 8'd3;
        rom[111][7] = -8'd1;
        rom[111][8] = 8'd8;
        rom[111][9] = 8'd13;
        rom[111][10] = -8'd22;
        rom[111][11] = -8'd7;
        rom[111][12] = 8'd7;
        rom[111][13] = -8'd5;
        rom[111][14] = -8'd10;
        rom[111][15] = -8'd8;
        rom[111][16] = -8'd4;
        rom[111][17] = 8'd7;
        rom[111][18] = 8'd19;
        rom[111][19] = -8'd10;
        rom[111][20] = 8'd5;
        rom[111][21] = 8'd10;
        rom[111][22] = -8'd31;
        rom[111][23] = -8'd5;
        rom[111][24] = 8'd22;
        rom[111][25] = -8'd4;
        rom[111][26] = -8'd6;
        rom[111][27] = -8'd19;
        rom[111][28] = -8'd20;
        rom[111][29] = -8'd3;
        rom[111][30] = -8'd8;
        rom[111][31] = -8'd88;
        rom[112][0] = 8'd6;
        rom[112][1] = -8'd67;
        rom[112][2] = 8'd7;
        rom[112][3] = -8'd16;
        rom[112][4] = -8'd41;
        rom[112][5] = 8'd26;
        rom[112][6] = 8'd3;
        rom[112][7] = 8'd8;
        rom[112][8] = -8'd5;
        rom[112][9] = 8'd12;
        rom[112][10] = -8'd4;
        rom[112][11] = -8'd29;
        rom[112][12] = -8'd19;
        rom[112][13] = 8'd6;
        rom[112][14] = -8'd19;
        rom[112][15] = 8'd26;
        rom[112][16] = -8'd59;
        rom[112][17] = 8'd26;
        rom[112][18] = 8'd17;
        rom[112][19] = -8'd16;
        rom[112][20] = 8'd10;
        rom[112][21] = 8'd4;
        rom[112][22] = -8'd33;
        rom[112][23] = 8'd1;
        rom[112][24] = -8'd55;
        rom[112][25] = -8'd8;
        rom[112][26] = -8'd3;
        rom[112][27] = -8'd3;
        rom[112][28] = 8'd29;
        rom[112][29] = 8'd9;
        rom[112][30] = -8'd45;
        rom[112][31] = 8'd8;
        rom[113][0] = -8'd19;
        rom[113][1] = -8'd1;
        rom[113][2] = -8'd2;
        rom[113][3] = -8'd4;
        rom[113][4] = 8'd44;
        rom[113][5] = 8'd24;
        rom[113][6] = -8'd24;
        rom[113][7] = -8'd20;
        rom[113][8] = -8'd33;
        rom[113][9] = 8'd7;
        rom[113][10] = 8'd1;
        rom[113][11] = 8'd20;
        rom[113][12] = 8'd1;
        rom[113][13] = 8'd46;
        rom[113][14] = -8'd31;
        rom[113][15] = -8'd32;
        rom[113][16] = 8'd9;
        rom[113][17] = 8'd7;
        rom[113][18] = -8'd17;
        rom[113][19] = 8'd11;
        rom[113][20] = -8'd22;
        rom[113][21] = 8'd21;
        rom[113][22] = -8'd21;
        rom[113][23] = -8'd17;
        rom[113][24] = 8'd5;
        rom[113][25] = 8'd6;
        rom[113][26] = 8'd3;
        rom[113][27] = -8'd6;
        rom[113][28] = 8'd17;
        rom[113][29] = 8'd6;
        rom[113][30] = -8'd14;
        rom[113][31] = 8'd10;
        rom[114][0] = -8'd16;
        rom[114][1] = 8'd14;
        rom[114][2] = -8'd31;
        rom[114][3] = 8'd3;
        rom[114][4] = 8'd13;
        rom[114][5] = 8'd9;
        rom[114][6] = -8'd5;
        rom[114][7] = -8'd1;
        rom[114][8] = 8'd19;
        rom[114][9] = -8'd16;
        rom[114][10] = -8'd13;
        rom[114][11] = -8'd6;
        rom[114][12] = 8'd19;
        rom[114][13] = 8'd10;
        rom[114][14] = 8'd9;
        rom[114][15] = -8'd26;
        rom[114][16] = 8'd20;
        rom[114][17] = -8'd3;
        rom[114][18] = -8'd20;
        rom[114][19] = 8'd10;
        rom[114][20] = 8'd2;
        rom[114][21] = 8'd2;
        rom[114][22] = -8'd25;
        rom[114][23] = 8'd0;
        rom[114][24] = -8'd1;
        rom[114][25] = -8'd1;
        rom[114][26] = -8'd14;
        rom[114][27] = -8'd17;
        rom[114][28] = -8'd14;
        rom[114][29] = -8'd8;
        rom[114][30] = -8'd19;
        rom[114][31] = -8'd20;
        rom[115][0] = 8'd22;
        rom[115][1] = -8'd26;
        rom[115][2] = 8'd19;
        rom[115][3] = 8'd2;
        rom[115][4] = 8'd22;
        rom[115][5] = 8'd8;
        rom[115][6] = -8'd4;
        rom[115][7] = -8'd27;
        rom[115][8] = 8'd16;
        rom[115][9] = 8'd16;
        rom[115][10] = 8'd7;
        rom[115][11] = 8'd8;
        rom[115][12] = 8'd0;
        rom[115][13] = 8'd23;
        rom[115][14] = -8'd5;
        rom[115][15] = -8'd29;
        rom[115][16] = -8'd1;
        rom[115][17] = 8'd31;
        rom[115][18] = -8'd19;
        rom[115][19] = 8'd8;
        rom[115][20] = 8'd4;
        rom[115][21] = -8'd12;
        rom[115][22] = 8'd51;
        rom[115][23] = -8'd18;
        rom[115][24] = 8'd2;
        rom[115][25] = 8'd5;
        rom[115][26] = -8'd59;
        rom[115][27] = 8'd1;
        rom[115][28] = -8'd15;
        rom[115][29] = -8'd23;
        rom[115][30] = 8'd10;
        rom[115][31] = -8'd5;
        rom[116][0] = 8'd16;
        rom[116][1] = -8'd59;
        rom[116][2] = -8'd18;
        rom[116][3] = 8'd48;
        rom[116][4] = -8'd7;
        rom[116][5] = -8'd17;
        rom[116][6] = -8'd20;
        rom[116][7] = -8'd3;
        rom[116][8] = 8'd6;
        rom[116][9] = 8'd16;
        rom[116][10] = -8'd4;
        rom[116][11] = -8'd7;
        rom[116][12] = -8'd15;
        rom[116][13] = 8'd18;
        rom[116][14] = 8'd14;
        rom[116][15] = -8'd21;
        rom[116][16] = -8'd23;
        rom[116][17] = 8'd38;
        rom[116][18] = -8'd5;
        rom[116][19] = -8'd10;
        rom[116][20] = -8'd51;
        rom[116][21] = -8'd6;
        rom[116][22] = 8'd7;
        rom[116][23] = -8'd21;
        rom[116][24] = -8'd38;
        rom[116][25] = -8'd22;
        rom[116][26] = 8'd16;
        rom[116][27] = -8'd13;
        rom[116][28] = -8'd35;
        rom[116][29] = -8'd45;
        rom[116][30] = -8'd38;
        rom[116][31] = -8'd3;
        rom[117][0] = 8'd31;
        rom[117][1] = -8'd3;
        rom[117][2] = -8'd53;
        rom[117][3] = 8'd31;
        rom[117][4] = 8'd6;
        rom[117][5] = 8'd9;
        rom[117][6] = 8'd22;
        rom[117][7] = 8'd23;
        rom[117][8] = -8'd7;
        rom[117][9] = -8'd61;
        rom[117][10] = 8'd1;
        rom[117][11] = 8'd8;
        rom[117][12] = 8'd16;
        rom[117][13] = -8'd14;
        rom[117][14] = 8'd26;
        rom[117][15] = -8'd25;
        rom[117][16] = 8'd12;
        rom[117][17] = 8'd6;
        rom[117][18] = -8'd28;
        rom[117][19] = -8'd33;
        rom[117][20] = 8'd24;
        rom[117][21] = 8'd28;
        rom[117][22] = 8'd30;
        rom[117][23] = -8'd11;
        rom[117][24] = 8'd17;
        rom[117][25] = 8'd5;
        rom[117][26] = -8'd4;
        rom[117][27] = -8'd11;
        rom[117][28] = -8'd11;
        rom[117][29] = 8'd4;
        rom[117][30] = 8'd7;
        rom[117][31] = -8'd128;
        rom[118][0] = 8'd12;
        rom[118][1] = -8'd40;
        rom[118][2] = -8'd26;
        rom[118][3] = 8'd20;
        rom[118][4] = -8'd4;
        rom[118][5] = 8'd9;
        rom[118][6] = -8'd11;
        rom[118][7] = -8'd14;
        rom[118][8] = 8'd15;
        rom[118][9] = 8'd22;
        rom[118][10] = -8'd11;
        rom[118][11] = 8'd10;
        rom[118][12] = -8'd1;
        rom[118][13] = 8'd13;
        rom[118][14] = -8'd4;
        rom[118][15] = -8'd4;
        rom[118][16] = -8'd52;
        rom[118][17] = 8'd18;
        rom[118][18] = 8'd22;
        rom[118][19] = -8'd3;
        rom[118][20] = 8'd24;
        rom[118][21] = 8'd2;
        rom[118][22] = -8'd27;
        rom[118][23] = -8'd5;
        rom[118][24] = -8'd14;
        rom[118][25] = -8'd33;
        rom[118][26] = 8'd3;
        rom[118][27] = 8'd12;
        rom[118][28] = 8'd0;
        rom[118][29] = -8'd4;
        rom[118][30] = 8'd10;
        rom[118][31] = 8'd5;
        rom[119][0] = 8'd20;
        rom[119][1] = 8'd15;
        rom[119][2] = -8'd30;
        rom[119][3] = -8'd2;
        rom[119][4] = 8'd9;
        rom[119][5] = 8'd3;
        rom[119][6] = 8'd40;
        rom[119][7] = 8'd36;
        rom[119][8] = -8'd9;
        rom[119][9] = -8'd42;
        rom[119][10] = 8'd28;
        rom[119][11] = 8'd12;
        rom[119][12] = 8'd0;
        rom[119][13] = -8'd12;
        rom[119][14] = 8'd15;
        rom[119][15] = -8'd15;
        rom[119][16] = -8'd7;
        rom[119][17] = 8'd3;
        rom[119][18] = -8'd9;
        rom[119][19] = -8'd1;
        rom[119][20] = 8'd30;
        rom[119][21] = 8'd21;
        rom[119][22] = 8'd5;
        rom[119][23] = 8'd9;
        rom[119][24] = 8'd3;
        rom[119][25] = 8'd10;
        rom[119][26] = -8'd13;
        rom[119][27] = 8'd12;
        rom[119][28] = -8'd15;
        rom[119][29] = 8'd25;
        rom[119][30] = 8'd18;
        rom[119][31] = -8'd62;
        rom[120][0] = 8'd13;
        rom[120][1] = -8'd37;
        rom[120][2] = -8'd3;
        rom[120][3] = -8'd24;
        rom[120][4] = -8'd21;
        rom[120][5] = -8'd25;
        rom[120][6] = 8'd29;
        rom[120][7] = 8'd6;
        rom[120][8] = -8'd9;
        rom[120][9] = -8'd23;
        rom[120][10] = 8'd0;
        rom[120][11] = -8'd18;
        rom[120][12] = -8'd4;
        rom[120][13] = -8'd4;
        rom[120][14] = -8'd2;
        rom[120][15] = 8'd5;
        rom[120][16] = -8'd35;
        rom[120][17] = 8'd19;
        rom[120][18] = 8'd5;
        rom[120][19] = -8'd53;
        rom[120][20] = -8'd47;
        rom[120][21] = -8'd15;
        rom[120][22] = 8'd0;
        rom[120][23] = 8'd23;
        rom[120][24] = -8'd34;
        rom[120][25] = -8'd10;
        rom[120][26] = 8'd50;
        rom[120][27] = 8'd19;
        rom[120][28] = 8'd12;
        rom[120][29] = -8'd18;
        rom[120][30] = -8'd15;
        rom[120][31] = -8'd4;
        rom[121][0] = 8'd8;
        rom[121][1] = -8'd12;
        rom[121][2] = -8'd15;
        rom[121][3] = -8'd51;
        rom[121][4] = 8'd2;
        rom[121][5] = 8'd12;
        rom[121][6] = -8'd18;
        rom[121][7] = -8'd8;
        rom[121][8] = -8'd81;
        rom[121][9] = 8'd11;
        rom[121][10] = 8'd14;
        rom[121][11] = -8'd18;
        rom[121][12] = -8'd23;
        rom[121][13] = -8'd9;
        rom[121][14] = 8'd2;
        rom[121][15] = 8'd4;
        rom[121][16] = -8'd12;
        rom[121][17] = 8'd29;
        rom[121][18] = 8'd9;
        rom[121][19] = -8'd37;
        rom[121][20] = -8'd20;
        rom[121][21] = -8'd25;
        rom[121][22] = 8'd8;
        rom[121][23] = -8'd18;
        rom[121][24] = 8'd13;
        rom[121][25] = 8'd24;
        rom[121][26] = 8'd14;
        rom[121][27] = 8'd18;
        rom[121][28] = -8'd1;
        rom[121][29] = -8'd21;
        rom[121][30] = -8'd17;
        rom[121][31] = -8'd5;
        rom[122][0] = 8'd12;
        rom[122][1] = -8'd7;
        rom[122][2] = -8'd45;
        rom[122][3] = 8'd17;
        rom[122][4] = -8'd31;
        rom[122][5] = 8'd2;
        rom[122][6] = -8'd13;
        rom[122][7] = -8'd11;
        rom[122][8] = -8'd29;
        rom[122][9] = 8'd19;
        rom[122][10] = -8'd8;
        rom[122][11] = 8'd36;
        rom[122][12] = 8'd27;
        rom[122][13] = 8'd11;
        rom[122][14] = 8'd44;
        rom[122][15] = -8'd21;
        rom[122][16] = -8'd10;
        rom[122][17] = 8'd7;
        rom[122][18] = 8'd1;
        rom[122][19] = 8'd32;
        rom[122][20] = -8'd18;
        rom[122][21] = -8'd23;
        rom[122][22] = 8'd8;
        rom[122][23] = -8'd4;
        rom[122][24] = -8'd8;
        rom[122][25] = -8'd11;
        rom[122][26] = 8'd16;
        rom[122][27] = 8'd10;
        rom[122][28] = -8'd3;
        rom[122][29] = 8'd15;
        rom[122][30] = -8'd53;
        rom[122][31] = -8'd20;
        rom[123][0] = 8'd10;
        rom[123][1] = 8'd11;
        rom[123][2] = -8'd69;
        rom[123][3] = 8'd26;
        rom[123][4] = -8'd13;
        rom[123][5] = 8'd11;
        rom[123][6] = 8'd4;
        rom[123][7] = 8'd11;
        rom[123][8] = 8'd19;
        rom[123][9] = -8'd4;
        rom[123][10] = -8'd8;
        rom[123][11] = 8'd24;
        rom[123][12] = -8'd3;
        rom[123][13] = 8'd10;
        rom[123][14] = 8'd8;
        rom[123][15] = -8'd12;
        rom[123][16] = 8'd11;
        rom[123][17] = -8'd19;
        rom[123][18] = -8'd43;
        rom[123][19] = -8'd50;
        rom[123][20] = 8'd23;
        rom[123][21] = 8'd44;
        rom[123][22] = 8'd8;
        rom[123][23] = -8'd39;
        rom[123][24] = 8'd36;
        rom[123][25] = 8'd9;
        rom[123][26] = -8'd3;
        rom[123][27] = 8'd4;
        rom[123][28] = -8'd8;
        rom[123][29] = -8'd6;
        rom[123][30] = 8'd33;
        rom[123][31] = -8'd74;
        rom[124][0] = 8'd3;
        rom[124][1] = 8'd10;
        rom[124][2] = 8'd8;
        rom[124][3] = -8'd9;
        rom[124][4] = -8'd18;
        rom[124][5] = -8'd19;
        rom[124][6] = 8'd10;
        rom[124][7] = -8'd2;
        rom[124][8] = 8'd32;
        rom[124][9] = -8'd30;
        rom[124][10] = 8'd6;
        rom[124][11] = -8'd19;
        rom[124][12] = -8'd25;
        rom[124][13] = -8'd7;
        rom[124][14] = -8'd2;
        rom[124][15] = 8'd9;
        rom[124][16] = 8'd55;
        rom[124][17] = -8'd22;
        rom[124][18] = -8'd3;
        rom[124][19] = -8'd24;
        rom[124][20] = -8'd2;
        rom[124][21] = -8'd10;
        rom[124][22] = 8'd2;
        rom[124][23] = -8'd33;
        rom[124][24] = 8'd0;
        rom[124][25] = -8'd30;
        rom[124][26] = -8'd9;
        rom[124][27] = -8'd1;
        rom[124][28] = -8'd27;
        rom[124][29] = 8'd19;
        rom[124][30] = -8'd22;
        rom[124][31] = -8'd7;
        rom[125][0] = -8'd10;
        rom[125][1] = 8'd21;
        rom[125][2] = 8'd22;
        rom[125][3] = 8'd20;
        rom[125][4] = 8'd13;
        rom[125][5] = 8'd1;
        rom[125][6] = 8'd21;
        rom[125][7] = 8'd7;
        rom[125][8] = -8'd22;
        rom[125][9] = 8'd30;
        rom[125][10] = 8'd23;
        rom[125][11] = 8'd30;
        rom[125][12] = 8'd1;
        rom[125][13] = 8'd10;
        rom[125][14] = 8'd35;
        rom[125][15] = 8'd4;
        rom[125][16] = 8'd11;
        rom[125][17] = -8'd14;
        rom[125][18] = 8'd14;
        rom[125][19] = -8'd5;
        rom[125][20] = 8'd9;
        rom[125][21] = 8'd6;
        rom[125][22] = -8'd9;
        rom[125][23] = 8'd28;
        rom[125][24] = 8'd5;
        rom[125][25] = 8'd15;
        rom[125][26] = -8'd9;
        rom[125][27] = 8'd3;
        rom[125][28] = -8'd40;
        rom[125][29] = 8'd5;
        rom[125][30] = -8'd22;
        rom[125][31] = -8'd26;
        rom[126][0] = 8'd37;
        rom[126][1] = -8'd7;
        rom[126][2] = -8'd41;
        rom[126][3] = -8'd23;
        rom[126][4] = 8'd16;
        rom[126][5] = 8'd16;
        rom[126][6] = -8'd22;
        rom[126][7] = -8'd2;
        rom[126][8] = 8'd17;
        rom[126][9] = 8'd18;
        rom[126][10] = -8'd18;
        rom[126][11] = 8'd16;
        rom[126][12] = 8'd14;
        rom[126][13] = 8'd38;
        rom[126][14] = 8'd15;
        rom[126][15] = -8'd4;
        rom[126][16] = -8'd16;
        rom[126][17] = -8'd7;
        rom[126][18] = -8'd57;
        rom[126][19] = -8'd2;
        rom[126][20] = 8'd17;
        rom[126][21] = 8'd37;
        rom[126][22] = 8'd16;
        rom[126][23] = -8'd19;
        rom[126][24] = -8'd14;
        rom[126][25] = 8'd2;
        rom[126][26] = 8'd27;
        rom[126][27] = 8'd3;
        rom[126][28] = 8'd17;
        rom[126][29] = 8'd51;
        rom[126][30] = 8'd26;
        rom[126][31] = -8'd17;
        rom[127][0] = -8'd6;
        rom[127][1] = 8'd17;
        rom[127][2] = -8'd82;
        rom[127][3] = 8'd16;
        rom[127][4] = 8'd25;
        rom[127][5] = 8'd18;
        rom[127][6] = -8'd5;
        rom[127][7] = 8'd19;
        rom[127][8] = 8'd4;
        rom[127][9] = -8'd3;
        rom[127][10] = -8'd9;
        rom[127][11] = 8'd20;
        rom[127][12] = 8'd18;
        rom[127][13] = -8'd27;
        rom[127][14] = 8'd7;
        rom[127][15] = 8'd0;
        rom[127][16] = 8'd20;
        rom[127][17] = 8'd8;
        rom[127][18] = -8'd9;
        rom[127][19] = 8'd5;
        rom[127][20] = 8'd13;
        rom[127][21] = 8'd44;
        rom[127][22] = -8'd11;
        rom[127][23] = -8'd37;
        rom[127][24] = 8'd27;
        rom[127][25] = -8'd15;
        rom[127][26] = -8'd8;
        rom[127][27] = 8'd27;
        rom[127][28] = -8'd25;
        rom[127][29] = 8'd11;
        rom[127][30] = 8'd17;
        rom[127][31] = -8'd78;
        rom[128][0] = -8'd16;
        rom[128][1] = -8'd26;
        rom[128][2] = 8'd17;
        rom[128][3] = -8'd4;
        rom[128][4] = -8'd2;
        rom[128][5] = 8'd43;
        rom[128][6] = -8'd32;
        rom[128][7] = 8'd0;
        rom[128][8] = -8'd14;
        rom[128][9] = -8'd6;
        rom[128][10] = -8'd40;
        rom[128][11] = 8'd18;
        rom[128][12] = 8'd19;
        rom[128][13] = -8'd2;
        rom[128][14] = -8'd16;
        rom[128][15] = -8'd5;
        rom[128][16] = -8'd9;
        rom[128][17] = 8'd9;
        rom[128][18] = 8'd3;
        rom[128][19] = 8'd15;
        rom[128][20] = 8'd17;
        rom[128][21] = 8'd19;
        rom[128][22] = -8'd34;
        rom[128][23] = -8'd13;
        rom[128][24] = -8'd40;
        rom[128][25] = -8'd12;
        rom[128][26] = -8'd16;
        rom[128][27] = -8'd29;
        rom[128][28] = 8'd28;
        rom[128][29] = 8'd8;
        rom[128][30] = -8'd57;
        rom[128][31] = 8'd9;
        rom[129][0] = -8'd19;
        rom[129][1] = -8'd6;
        rom[129][2] = -8'd13;
        rom[129][3] = -8'd9;
        rom[129][4] = -8'd25;
        rom[129][5] = 8'd3;
        rom[129][6] = 8'd48;
        rom[129][7] = 8'd17;
        rom[129][8] = -8'd25;
        rom[129][9] = -8'd19;
        rom[129][10] = 8'd26;
        rom[129][11] = 8'd48;
        rom[129][12] = -8'd9;
        rom[129][13] = 8'd17;
        rom[129][14] = -8'd30;
        rom[129][15] = 8'd24;
        rom[129][16] = -8'd23;
        rom[129][17] = 8'd9;
        rom[129][18] = 8'd8;
        rom[129][19] = -8'd3;
        rom[129][20] = 8'd32;
        rom[129][21] = 8'd15;
        rom[129][22] = -8'd18;
        rom[129][23] = 8'd15;
        rom[129][24] = -8'd1;
        rom[129][25] = -8'd34;
        rom[129][26] = 8'd17;
        rom[129][27] = 8'd15;
        rom[129][28] = -8'd10;
        rom[129][29] = 8'd39;
        rom[129][30] = 8'd0;
        rom[129][31] = 8'd15;
        rom[130][0] = -8'd32;
        rom[130][1] = 8'd1;
        rom[130][2] = 8'd7;
        rom[130][3] = 8'd18;
        rom[130][4] = -8'd9;
        rom[130][5] = -8'd4;
        rom[130][6] = 8'd7;
        rom[130][7] = 8'd10;
        rom[130][8] = -8'd13;
        rom[130][9] = -8'd37;
        rom[130][10] = -8'd6;
        rom[130][11] = -8'd12;
        rom[130][12] = 8'd3;
        rom[130][13] = 8'd9;
        rom[130][14] = -8'd34;
        rom[130][15] = -8'd25;
        rom[130][16] = 8'd12;
        rom[130][17] = 8'd8;
        rom[130][18] = -8'd2;
        rom[130][19] = 8'd28;
        rom[130][20] = -8'd6;
        rom[130][21] = -8'd16;
        rom[130][22] = -8'd7;
        rom[130][23] = -8'd59;
        rom[130][24] = -8'd20;
        rom[130][25] = -8'd6;
        rom[130][26] = -8'd22;
        rom[130][27] = -8'd12;
        rom[130][28] = 8'd26;
        rom[130][29] = -8'd28;
        rom[130][30] = 8'd11;
        rom[130][31] = 8'd21;
        rom[131][0] = -8'd12;
        rom[131][1] = -8'd67;
        rom[131][2] = -8'd12;
        rom[131][3] = -8'd25;
        rom[131][4] = -8'd14;
        rom[131][5] = -8'd4;
        rom[131][6] = 8'd42;
        rom[131][7] = 8'd1;
        rom[131][8] = -8'd21;
        rom[131][9] = 8'd9;
        rom[131][10] = 8'd12;
        rom[131][11] = 8'd40;
        rom[131][12] = 8'd32;
        rom[131][13] = 8'd20;
        rom[131][14] = -8'd41;
        rom[131][15] = -8'd33;
        rom[131][16] = -8'd1;
        rom[131][17] = 8'd4;
        rom[131][18] = -8'd37;
        rom[131][19] = -8'd7;
        rom[131][20] = 8'd24;
        rom[131][21] = 8'd3;
        rom[131][22] = 8'd47;
        rom[131][23] = -8'd2;
        rom[131][24] = -8'd3;
        rom[131][25] = -8'd29;
        rom[131][26] = -8'd8;
        rom[131][27] = -8'd5;
        rom[131][28] = -8'd3;
        rom[131][29] = 8'd10;
        rom[131][30] = -8'd11;
        rom[131][31] = 8'd14;
        rom[132][0] = -8'd7;
        rom[132][1] = -8'd65;
        rom[132][2] = -8'd22;
        rom[132][3] = 8'd31;
        rom[132][4] = 8'd27;
        rom[132][5] = 8'd21;
        rom[132][6] = -8'd13;
        rom[132][7] = 8'd8;
        rom[132][8] = 8'd3;
        rom[132][9] = 8'd13;
        rom[132][10] = -8'd7;
        rom[132][11] = 8'd27;
        rom[132][12] = -8'd13;
        rom[132][13] = 8'd33;
        rom[132][14] = -8'd3;
        rom[132][15] = -8'd14;
        rom[132][16] = -8'd24;
        rom[132][17] = 8'd28;
        rom[132][18] = 8'd13;
        rom[132][19] = -8'd19;
        rom[132][20] = -8'd18;
        rom[132][21] = 8'd46;
        rom[132][22] = -8'd2;
        rom[132][23] = 8'd3;
        rom[132][24] = -8'd10;
        rom[132][25] = -8'd16;
        rom[132][26] = -8'd14;
        rom[132][27] = -8'd2;
        rom[132][28] = -8'd5;
        rom[132][29] = -8'd18;
        rom[132][30] = -8'd36;
        rom[132][31] = 8'd19;
        rom[133][0] = -8'd1;
        rom[133][1] = -8'd14;
        rom[133][2] = 8'd16;
        rom[133][3] = 8'd27;
        rom[133][4] = -8'd29;
        rom[133][5] = 8'd8;
        rom[133][6] = 8'd16;
        rom[133][7] = 8'd11;
        rom[133][8] = -8'd19;
        rom[133][9] = -8'd35;
        rom[133][10] = 8'd22;
        rom[133][11] = 8'd10;
        rom[133][12] = -8'd11;
        rom[133][13] = 8'd19;
        rom[133][14] = 8'd0;
        rom[133][15] = -8'd19;
        rom[133][16] = 8'd24;
        rom[133][17] = -8'd34;
        rom[133][18] = 8'd7;
        rom[133][19] = -8'd30;
        rom[133][20] = -8'd4;
        rom[133][21] = 8'd4;
        rom[133][22] = 8'd28;
        rom[133][23] = -8'd14;
        rom[133][24] = 8'd7;
        rom[133][25] = 8'd54;
        rom[133][26] = 8'd10;
        rom[133][27] = -8'd15;
        rom[133][28] = 8'd27;
        rom[133][29] = -8'd10;
        rom[133][30] = -8'd11;
        rom[133][31] = -8'd51;
        rom[134][0] = 8'd17;
        rom[134][1] = -8'd19;
        rom[134][2] = -8'd22;
        rom[134][3] = -8'd12;
        rom[134][4] = 8'd26;
        rom[134][5] = -8'd16;
        rom[134][6] = -8'd6;
        rom[134][7] = 8'd2;
        rom[134][8] = -8'd20;
        rom[134][9] = 8'd17;
        rom[134][10] = -8'd1;
        rom[134][11] = 8'd18;
        rom[134][12] = 8'd15;
        rom[134][13] = 8'd2;
        rom[134][14] = 8'd18;
        rom[134][15] = -8'd1;
        rom[134][16] = -8'd48;
        rom[134][17] = 8'd22;
        rom[134][18] = 8'd15;
        rom[134][19] = 8'd11;
        rom[134][20] = 8'd13;
        rom[134][21] = 8'd11;
        rom[134][22] = -8'd10;
        rom[134][23] = 8'd13;
        rom[134][24] = 8'd6;
        rom[134][25] = -8'd32;
        rom[134][26] = -8'd19;
        rom[134][27] = 8'd25;
        rom[134][28] = -8'd3;
        rom[134][29] = 8'd4;
        rom[134][30] = 8'd24;
        rom[134][31] = 8'd53;
        rom[135][0] = 8'd25;
        rom[135][1] = -8'd5;
        rom[135][2] = 8'd11;
        rom[135][3] = -8'd4;
        rom[135][4] = -8'd13;
        rom[135][5] = -8'd2;
        rom[135][6] = 8'd11;
        rom[135][7] = 8'd21;
        rom[135][8] = 8'd11;
        rom[135][9] = -8'd18;
        rom[135][10] = 8'd36;
        rom[135][11] = -8'd20;
        rom[135][12] = -8'd23;
        rom[135][13] = -8'd32;
        rom[135][14] = -8'd9;
        rom[135][15] = 8'd13;
        rom[135][16] = 8'd31;
        rom[135][17] = -8'd4;
        rom[135][18] = 8'd34;
        rom[135][19] = -8'd2;
        rom[135][20] = 8'd23;
        rom[135][21] = -8'd49;
        rom[135][22] = 8'd2;
        rom[135][23] = 8'd2;
        rom[135][24] = 8'd33;
        rom[135][25] = 8'd13;
        rom[135][26] = 8'd0;
        rom[135][27] = 8'd21;
        rom[135][28] = 8'd9;
        rom[135][29] = 8'd2;
        rom[135][30] = -8'd4;
        rom[135][31] = -8'd10;
        rom[136][0] = 8'd8;
        rom[136][1] = -8'd9;
        rom[136][2] = 8'd25;
        rom[136][3] = -8'd9;
        rom[136][4] = -8'd10;
        rom[136][5] = 8'd16;
        rom[136][6] = 8'd3;
        rom[136][7] = 8'd18;
        rom[136][8] = 8'd5;
        rom[136][9] = -8'd22;
        rom[136][10] = 8'd4;
        rom[136][11] = 8'd10;
        rom[136][12] = 8'd6;
        rom[136][13] = -8'd4;
        rom[136][14] = -8'd3;
        rom[136][15] = 8'd11;
        rom[136][16] = -8'd27;
        rom[136][17] = 8'd4;
        rom[136][18] = 8'd12;
        rom[136][19] = -8'd59;
        rom[136][20] = -8'd7;
        rom[136][21] = 8'd17;
        rom[136][22] = -8'd1;
        rom[136][23] = 8'd24;
        rom[136][24] = 8'd4;
        rom[136][25] = -8'd1;
        rom[136][26] = 8'd44;
        rom[136][27] = 8'd2;
        rom[136][28] = 8'd17;
        rom[136][29] = 8'd3;
        rom[136][30] = -8'd45;
        rom[136][31] = 8'd14;
        rom[137][0] = 8'd7;
        rom[137][1] = 8'd33;
        rom[137][2] = 8'd0;
        rom[137][3] = -8'd38;
        rom[137][4] = -8'd7;
        rom[137][5] = 8'd28;
        rom[137][6] = -8'd27;
        rom[137][7] = 8'd4;
        rom[137][8] = -8'd87;
        rom[137][9] = 8'd28;
        rom[137][10] = 8'd11;
        rom[137][11] = 8'd12;
        rom[137][12] = 8'd19;
        rom[137][13] = 8'd1;
        rom[137][14] = -8'd24;
        rom[137][15] = 8'd12;
        rom[137][16] = 8'd1;
        rom[137][17] = 8'd3;
        rom[137][18] = 8'd16;
        rom[137][19] = 8'd1;
        rom[137][20] = -8'd18;
        rom[137][21] = 8'd7;
        rom[137][22] = -8'd33;
        rom[137][23] = -8'd7;
        rom[137][24] = 8'd23;
        rom[137][25] = -8'd8;
        rom[137][26] = 8'd26;
        rom[137][27] = -8'd6;
        rom[137][28] = 8'd18;
        rom[137][29] = -8'd8;
        rom[137][30] = -8'd28;
        rom[137][31] = 8'd1;
        rom[138][0] = 8'd8;
        rom[138][1] = -8'd27;
        rom[138][2] = -8'd13;
        rom[138][3] = 8'd3;
        rom[138][4] = -8'd15;
        rom[138][5] = -8'd38;
        rom[138][6] = -8'd9;
        rom[138][7] = -8'd6;
        rom[138][8] = -8'd20;
        rom[138][9] = -8'd23;
        rom[138][10] = -8'd13;
        rom[138][11] = -8'd3;
        rom[138][12] = 8'd2;
        rom[138][13] = 8'd20;
        rom[138][14] = 8'd19;
        rom[138][15] = 8'd13;
        rom[138][16] = -8'd1;
        rom[138][17] = -8'd11;
        rom[138][18] = 8'd26;
        rom[138][19] = 8'd36;
        rom[138][20] = 8'd1;
        rom[138][21] = -8'd21;
        rom[138][22] = 8'd17;
        rom[138][23] = -8'd30;
        rom[138][24] = -8'd12;
        rom[138][25] = -8'd51;
        rom[138][26] = 8'd26;
        rom[138][27] = 8'd8;
        rom[138][28] = -8'd2;
        rom[138][29] = 8'd12;
        rom[138][30] = -8'd9;
        rom[138][31] = -8'd7;
        rom[139][0] = -8'd5;
        rom[139][1] = 8'd7;
        rom[139][2] = -8'd3;
        rom[139][3] = 8'd23;
        rom[139][4] = -8'd44;
        rom[139][5] = -8'd8;
        rom[139][6] = -8'd2;
        rom[139][7] = 8'd8;
        rom[139][8] = 8'd21;
        rom[139][9] = -8'd2;
        rom[139][10] = 8'd5;
        rom[139][11] = 8'd11;
        rom[139][12] = -8'd8;
        rom[139][13] = 8'd46;
        rom[139][14] = 8'd26;
        rom[139][15] = 8'd37;
        rom[139][16] = 8'd5;
        rom[139][17] = -8'd27;
        rom[139][18] = -8'd6;
        rom[139][19] = 8'd0;
        rom[139][20] = 8'd21;
        rom[139][21] = -8'd18;
        rom[139][22] = -8'd5;
        rom[139][23] = -8'd56;
        rom[139][24] = 8'd21;
        rom[139][25] = -8'd36;
        rom[139][26] = 8'd1;
        rom[139][27] = -8'd7;
        rom[139][28] = 8'd33;
        rom[139][29] = -8'd6;
        rom[139][30] = 8'd12;
        rom[139][31] = 8'd4;
        rom[140][0] = 8'd4;
        rom[140][1] = -8'd28;
        rom[140][2] = 8'd36;
        rom[140][3] = 8'd4;
        rom[140][4] = 8'd25;
        rom[140][5] = 8'd2;
        rom[140][6] = 8'd34;
        rom[140][7] = -8'd7;
        rom[140][8] = -8'd12;
        rom[140][9] = 8'd0;
        rom[140][10] = 8'd13;
        rom[140][11] = -8'd2;
        rom[140][12] = -8'd48;
        rom[140][13] = 8'd2;
        rom[140][14] = -8'd15;
        rom[140][15] = -8'd9;
        rom[140][16] = 8'd50;
        rom[140][17] = -8'd14;
        rom[140][18] = 8'd11;
        rom[140][19] = -8'd17;
        rom[140][20] = -8'd22;
        rom[140][21] = 8'd3;
        rom[140][22] = -8'd7;
        rom[140][23] = -8'd20;
        rom[140][24] = 8'd0;
        rom[140][25] = 8'd9;
        rom[140][26] = -8'd3;
        rom[140][27] = -8'd2;
        rom[140][28] = -8'd16;
        rom[140][29] = 8'd4;
        rom[140][30] = -8'd62;
        rom[140][31] = 8'd0;
        rom[141][0] = -8'd12;
        rom[141][1] = -8'd7;
        rom[141][2] = 8'd38;
        rom[141][3] = -8'd12;
        rom[141][4] = 8'd22;
        rom[141][5] = -8'd7;
        rom[141][6] = -8'd7;
        rom[141][7] = -8'd40;
        rom[141][8] = -8'd13;
        rom[141][9] = 8'd10;
        rom[141][10] = 8'd17;
        rom[141][11] = -8'd3;
        rom[141][12] = -8'd15;
        rom[141][13] = -8'd5;
        rom[141][14] = 8'd24;
        rom[141][15] = -8'd27;
        rom[141][16] = 8'd3;
        rom[141][17] = 8'd0;
        rom[141][18] = 8'd31;
        rom[141][19] = 8'd24;
        rom[141][20] = -8'd31;
        rom[141][21] = -8'd34;
        rom[141][22] = 8'd4;
        rom[141][23] = -8'd3;
        rom[141][24] = 8'd6;
        rom[141][25] = 8'd28;
        rom[141][26] = -8'd11;
        rom[141][27] = -8'd28;
        rom[141][28] = -8'd13;
        rom[141][29] = -8'd36;
        rom[141][30] = -8'd5;
        rom[141][31] = 8'd6;
        rom[142][0] = 8'd40;
        rom[142][1] = 8'd32;
        rom[142][2] = -8'd56;
        rom[142][3] = -8'd23;
        rom[142][4] = -8'd12;
        rom[142][5] = -8'd30;
        rom[142][6] = -8'd55;
        rom[142][7] = 8'd5;
        rom[142][8] = 8'd15;
        rom[142][9] = -8'd17;
        rom[142][10] = 8'd25;
        rom[142][11] = 8'd26;
        rom[142][12] = -8'd9;
        rom[142][13] = -8'd23;
        rom[142][14] = 8'd9;
        rom[142][15] = -8'd15;
        rom[142][16] = 8'd5;
        rom[142][17] = -8'd43;
        rom[142][18] = -8'd19;
        rom[142][19] = 8'd20;
        rom[142][20] = 8'd11;
        rom[142][21] = 8'd0;
        rom[142][22] = 8'd29;
        rom[142][23] = -8'd12;
        rom[142][24] = -8'd16;
        rom[142][25] = -8'd9;
        rom[142][26] = 8'd12;
        rom[142][27] = -8'd31;
        rom[142][28] = -8'd2;
        rom[142][29] = 8'd23;
        rom[142][30] = 8'd1;
        rom[142][31] = 8'd0;
        rom[143][0] = 8'd11;
        rom[143][1] = -8'd18;
        rom[143][2] = -8'd35;
        rom[143][3] = 8'd0;
        rom[143][4] = 8'd24;
        rom[143][5] = -8'd2;
        rom[143][6] = 8'd8;
        rom[143][7] = 8'd17;
        rom[143][8] = 8'd1;
        rom[143][9] = 8'd18;
        rom[143][10] = 8'd8;
        rom[143][11] = -8'd5;
        rom[143][12] = 8'd4;
        rom[143][13] = -8'd28;
        rom[143][14] = 8'd31;
        rom[143][15] = -8'd3;
        rom[143][16] = 8'd20;
        rom[143][17] = 8'd21;
        rom[143][18] = 8'd15;
        rom[143][19] = 8'd21;
        rom[143][20] = -8'd1;
        rom[143][21] = -8'd16;
        rom[143][22] = 8'd2;
        rom[143][23] = -8'd11;
        rom[143][24] = 8'd21;
        rom[143][25] = -8'd1;
        rom[143][26] = 8'd11;
        rom[143][27] = -8'd17;
        rom[143][28] = 8'd15;
        rom[143][29] = 8'd17;
        rom[143][30] = 8'd36;
        rom[143][31] = -8'd6;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
