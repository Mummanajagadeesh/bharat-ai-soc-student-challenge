module rom_04_conv2d_3_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:287][0:31];

    initial begin
        rom[0][0] = 8'd16;
        rom[0][1] = -8'd2;
        rom[0][2] = 8'd23;
        rom[0][3] = -8'd42;
        rom[0][4] = 8'd23;
        rom[0][5] = -8'd40;
        rom[0][6] = 8'd20;
        rom[0][7] = 8'd4;
        rom[0][8] = -8'd3;
        rom[0][9] = 8'd18;
        rom[0][10] = 8'd19;
        rom[0][11] = -8'd17;
        rom[0][12] = -8'd4;
        rom[0][13] = -8'd29;
        rom[0][14] = 8'd1;
        rom[0][15] = -8'd30;
        rom[0][16] = -8'd10;
        rom[0][17] = 8'd5;
        rom[0][18] = -8'd12;
        rom[0][19] = 8'd7;
        rom[0][20] = 8'd0;
        rom[0][21] = 8'd10;
        rom[0][22] = -8'd3;
        rom[0][23] = -8'd1;
        rom[0][24] = 8'd13;
        rom[0][25] = 8'd24;
        rom[0][26] = -8'd2;
        rom[0][27] = 8'd13;
        rom[0][28] = -8'd8;
        rom[0][29] = -8'd9;
        rom[0][30] = 8'd2;
        rom[0][31] = 8'd4;
        rom[1][0] = 8'd40;
        rom[1][1] = 8'd22;
        rom[1][2] = -8'd32;
        rom[1][3] = 8'd3;
        rom[1][4] = -8'd18;
        rom[1][5] = 8'd16;
        rom[1][6] = -8'd26;
        rom[1][7] = -8'd63;
        rom[1][8] = -8'd10;
        rom[1][9] = -8'd8;
        rom[1][10] = 8'd8;
        rom[1][11] = -8'd1;
        rom[1][12] = -8'd16;
        rom[1][13] = 8'd18;
        rom[1][14] = 8'd3;
        rom[1][15] = 8'd0;
        rom[1][16] = 8'd20;
        rom[1][17] = 8'd15;
        rom[1][18] = -8'd1;
        rom[1][19] = 8'd5;
        rom[1][20] = 8'd8;
        rom[1][21] = 8'd10;
        rom[1][22] = 8'd25;
        rom[1][23] = 8'd15;
        rom[1][24] = 8'd8;
        rom[1][25] = -8'd18;
        rom[1][26] = 8'd12;
        rom[1][27] = -8'd12;
        rom[1][28] = 8'd1;
        rom[1][29] = -8'd3;
        rom[1][30] = -8'd35;
        rom[1][31] = 8'd24;
        rom[2][0] = -8'd34;
        rom[2][1] = 8'd21;
        rom[2][2] = 8'd5;
        rom[2][3] = -8'd36;
        rom[2][4] = 8'd2;
        rom[2][5] = 8'd28;
        rom[2][6] = -8'd6;
        rom[2][7] = 8'd4;
        rom[2][8] = 8'd67;
        rom[2][9] = -8'd61;
        rom[2][10] = -8'd32;
        rom[2][11] = 8'd16;
        rom[2][12] = -8'd7;
        rom[2][13] = -8'd17;
        rom[2][14] = -8'd10;
        rom[2][15] = -8'd18;
        rom[2][16] = 8'd31;
        rom[2][17] = 8'd19;
        rom[2][18] = -8'd27;
        rom[2][19] = -8'd9;
        rom[2][20] = -8'd26;
        rom[2][21] = -8'd29;
        rom[2][22] = 8'd15;
        rom[2][23] = -8'd41;
        rom[2][24] = -8'd39;
        rom[2][25] = 8'd42;
        rom[2][26] = -8'd33;
        rom[2][27] = -8'd26;
        rom[2][28] = 8'd8;
        rom[2][29] = -8'd7;
        rom[2][30] = -8'd18;
        rom[2][31] = 8'd21;
        rom[3][0] = 8'd37;
        rom[3][1] = -8'd29;
        rom[3][2] = -8'd5;
        rom[3][3] = 8'd0;
        rom[3][4] = 8'd2;
        rom[3][5] = -8'd12;
        rom[3][6] = -8'd7;
        rom[3][7] = -8'd27;
        rom[3][8] = 8'd30;
        rom[3][9] = 8'd16;
        rom[3][10] = 8'd2;
        rom[3][11] = 8'd29;
        rom[3][12] = -8'd15;
        rom[3][13] = 8'd14;
        rom[3][14] = 8'd2;
        rom[3][15] = -8'd63;
        rom[3][16] = 8'd24;
        rom[3][17] = -8'd1;
        rom[3][18] = -8'd6;
        rom[3][19] = 8'd14;
        rom[3][20] = -8'd13;
        rom[3][21] = 8'd1;
        rom[3][22] = -8'd3;
        rom[3][23] = -8'd29;
        rom[3][24] = -8'd7;
        rom[3][25] = -8'd23;
        rom[3][26] = -8'd15;
        rom[3][27] = 8'd9;
        rom[3][28] = -8'd23;
        rom[3][29] = 8'd5;
        rom[3][30] = 8'd13;
        rom[3][31] = 8'd32;
        rom[4][0] = -8'd36;
        rom[4][1] = 8'd2;
        rom[4][2] = -8'd1;
        rom[4][3] = 8'd58;
        rom[4][4] = -8'd15;
        rom[4][5] = -8'd12;
        rom[4][6] = 8'd27;
        rom[4][7] = -8'd28;
        rom[4][8] = -8'd32;
        rom[4][9] = -8'd8;
        rom[4][10] = -8'd8;
        rom[4][11] = 8'd32;
        rom[4][12] = 8'd12;
        rom[4][13] = -8'd19;
        rom[4][14] = -8'd14;
        rom[4][15] = 8'd27;
        rom[4][16] = -8'd8;
        rom[4][17] = 8'd40;
        rom[4][18] = 8'd24;
        rom[4][19] = -8'd44;
        rom[4][20] = 8'd13;
        rom[4][21] = -8'd17;
        rom[4][22] = -8'd22;
        rom[4][23] = 8'd13;
        rom[4][24] = 8'd28;
        rom[4][25] = -8'd11;
        rom[4][26] = -8'd32;
        rom[4][27] = -8'd17;
        rom[4][28] = -8'd7;
        rom[4][29] = -8'd8;
        rom[4][30] = -8'd18;
        rom[4][31] = 8'd1;
        rom[5][0] = -8'd1;
        rom[5][1] = 8'd34;
        rom[5][2] = -8'd7;
        rom[5][3] = -8'd12;
        rom[5][4] = -8'd19;
        rom[5][5] = -8'd3;
        rom[5][6] = -8'd14;
        rom[5][7] = 8'd20;
        rom[5][8] = 8'd11;
        rom[5][9] = -8'd8;
        rom[5][10] = 8'd36;
        rom[5][11] = 8'd10;
        rom[5][12] = -8'd13;
        rom[5][13] = 8'd30;
        rom[5][14] = 8'd25;
        rom[5][15] = -8'd68;
        rom[5][16] = -8'd17;
        rom[5][17] = 8'd2;
        rom[5][18] = -8'd43;
        rom[5][19] = -8'd16;
        rom[5][20] = -8'd2;
        rom[5][21] = 8'd4;
        rom[5][22] = -8'd15;
        rom[5][23] = -8'd49;
        rom[5][24] = -8'd31;
        rom[5][25] = 8'd28;
        rom[5][26] = -8'd45;
        rom[5][27] = -8'd2;
        rom[5][28] = 8'd9;
        rom[5][29] = -8'd7;
        rom[5][30] = 8'd20;
        rom[5][31] = 8'd47;
        rom[6][0] = -8'd7;
        rom[6][1] = 8'd26;
        rom[6][2] = -8'd35;
        rom[6][3] = -8'd22;
        rom[6][4] = -8'd23;
        rom[6][5] = -8'd23;
        rom[6][6] = -8'd26;
        rom[6][7] = 8'd1;
        rom[6][8] = 8'd19;
        rom[6][9] = -8'd27;
        rom[6][10] = 8'd13;
        rom[6][11] = 8'd17;
        rom[6][12] = 8'd16;
        rom[6][13] = 8'd20;
        rom[6][14] = 8'd29;
        rom[6][15] = 8'd42;
        rom[6][16] = -8'd16;
        rom[6][17] = -8'd21;
        rom[6][18] = -8'd38;
        rom[6][19] = 8'd2;
        rom[6][20] = 8'd28;
        rom[6][21] = 8'd19;
        rom[6][22] = 8'd19;
        rom[6][23] = 8'd0;
        rom[6][24] = 8'd14;
        rom[6][25] = -8'd6;
        rom[6][26] = -8'd8;
        rom[6][27] = -8'd34;
        rom[6][28] = 8'd20;
        rom[6][29] = -8'd5;
        rom[6][30] = -8'd7;
        rom[6][31] = 8'd16;
        rom[7][0] = 8'd2;
        rom[7][1] = -8'd7;
        rom[7][2] = 8'd3;
        rom[7][3] = 8'd5;
        rom[7][4] = 8'd7;
        rom[7][5] = -8'd35;
        rom[7][6] = 8'd2;
        rom[7][7] = 8'd1;
        rom[7][8] = -8'd59;
        rom[7][9] = 8'd15;
        rom[7][10] = 8'd11;
        rom[7][11] = 8'd1;
        rom[7][12] = -8'd2;
        rom[7][13] = 8'd17;
        rom[7][14] = -8'd19;
        rom[7][15] = -8'd7;
        rom[7][16] = -8'd4;
        rom[7][17] = 8'd2;
        rom[7][18] = 8'd7;
        rom[7][19] = 8'd3;
        rom[7][20] = 8'd2;
        rom[7][21] = 8'd10;
        rom[7][22] = 8'd11;
        rom[7][23] = 8'd14;
        rom[7][24] = -8'd15;
        rom[7][25] = 8'd7;
        rom[7][26] = 8'd26;
        rom[7][27] = 8'd16;
        rom[7][28] = -8'd8;
        rom[7][29] = 8'd5;
        rom[7][30] = -8'd6;
        rom[7][31] = 8'd9;
        rom[8][0] = 8'd13;
        rom[8][1] = -8'd4;
        rom[8][2] = 8'd8;
        rom[8][3] = 8'd28;
        rom[8][4] = 8'd14;
        rom[8][5] = 8'd26;
        rom[8][6] = -8'd6;
        rom[8][7] = 8'd29;
        rom[8][8] = -8'd54;
        rom[8][9] = 8'd36;
        rom[8][10] = 8'd34;
        rom[8][11] = 8'd8;
        rom[8][12] = -8'd17;
        rom[8][13] = 8'd18;
        rom[8][14] = 8'd7;
        rom[8][15] = -8'd13;
        rom[8][16] = 8'd24;
        rom[8][17] = 8'd6;
        rom[8][18] = -8'd2;
        rom[8][19] = -8'd6;
        rom[8][20] = 8'd38;
        rom[8][21] = 8'd21;
        rom[8][22] = 8'd18;
        rom[8][23] = 8'd9;
        rom[8][24] = -8'd11;
        rom[8][25] = -8'd22;
        rom[8][26] = 8'd13;
        rom[8][27] = 8'd36;
        rom[8][28] = -8'd3;
        rom[8][29] = 8'd12;
        rom[8][30] = 8'd20;
        rom[8][31] = -8'd64;
        rom[9][0] = -8'd1;
        rom[9][1] = 8'd13;
        rom[9][2] = -8'd24;
        rom[9][3] = -8'd18;
        rom[9][4] = 8'd24;
        rom[9][5] = 8'd3;
        rom[9][6] = -8'd9;
        rom[9][7] = 8'd46;
        rom[9][8] = 8'd75;
        rom[9][9] = 8'd15;
        rom[9][10] = 8'd18;
        rom[9][11] = -8'd12;
        rom[9][12] = -8'd21;
        rom[9][13] = -8'd1;
        rom[9][14] = 8'd13;
        rom[9][15] = 8'd23;
        rom[9][16] = -8'd1;
        rom[9][17] = 8'd16;
        rom[9][18] = -8'd5;
        rom[9][19] = 8'd4;
        rom[9][20] = -8'd6;
        rom[9][21] = -8'd1;
        rom[9][22] = 8'd20;
        rom[9][23] = -8'd21;
        rom[9][24] = 8'd27;
        rom[9][25] = 8'd11;
        rom[9][26] = 8'd2;
        rom[9][27] = -8'd29;
        rom[9][28] = -8'd1;
        rom[9][29] = 8'd9;
        rom[9][30] = 8'd27;
        rom[9][31] = 8'd0;
        rom[10][0] = -8'd29;
        rom[10][1] = 8'd10;
        rom[10][2] = -8'd8;
        rom[10][3] = -8'd40;
        rom[10][4] = -8'd19;
        rom[10][5] = 8'd7;
        rom[10][6] = 8'd9;
        rom[10][7] = 8'd54;
        rom[10][8] = -8'd22;
        rom[10][9] = 8'd42;
        rom[10][10] = -8'd9;
        rom[10][11] = 8'd24;
        rom[10][12] = 8'd32;
        rom[10][13] = -8'd46;
        rom[10][14] = -8'd6;
        rom[10][15] = 8'd30;
        rom[10][16] = -8'd1;
        rom[10][17] = 8'd13;
        rom[10][18] = -8'd41;
        rom[10][19] = -8'd10;
        rom[10][20] = 8'd25;
        rom[10][21] = 8'd39;
        rom[10][22] = 8'd10;
        rom[10][23] = -8'd8;
        rom[10][24] = 8'd39;
        rom[10][25] = 8'd10;
        rom[10][26] = 8'd21;
        rom[10][27] = 8'd9;
        rom[10][28] = 8'd10;
        rom[10][29] = 8'd2;
        rom[10][30] = 8'd44;
        rom[10][31] = -8'd10;
        rom[11][0] = 8'd6;
        rom[11][1] = -8'd14;
        rom[11][2] = -8'd2;
        rom[11][3] = 8'd2;
        rom[11][4] = -8'd15;
        rom[11][5] = -8'd29;
        rom[11][6] = 8'd9;
        rom[11][7] = 8'd25;
        rom[11][8] = -8'd53;
        rom[11][9] = -8'd16;
        rom[11][10] = -8'd2;
        rom[11][11] = -8'd12;
        rom[11][12] = 8'd34;
        rom[11][13] = -8'd17;
        rom[11][14] = -8'd28;
        rom[11][15] = 8'd4;
        rom[11][16] = -8'd51;
        rom[11][17] = -8'd18;
        rom[11][18] = 8'd21;
        rom[11][19] = -8'd10;
        rom[11][20] = -8'd3;
        rom[11][21] = 8'd21;
        rom[11][22] = -8'd10;
        rom[11][23] = 8'd7;
        rom[11][24] = 8'd0;
        rom[11][25] = -8'd3;
        rom[11][26] = -8'd6;
        rom[11][27] = 8'd12;
        rom[11][28] = -8'd4;
        rom[11][29] = -8'd17;
        rom[11][30] = 8'd16;
        rom[11][31] = 8'd33;
        rom[12][0] = 8'd35;
        rom[12][1] = 8'd36;
        rom[12][2] = 8'd10;
        rom[12][3] = -8'd7;
        rom[12][4] = -8'd1;
        rom[12][5] = 8'd4;
        rom[12][6] = -8'd2;
        rom[12][7] = 8'd23;
        rom[12][8] = 8'd23;
        rom[12][9] = -8'd18;
        rom[12][10] = 8'd27;
        rom[12][11] = -8'd27;
        rom[12][12] = -8'd29;
        rom[12][13] = 8'd18;
        rom[12][14] = 8'd12;
        rom[12][15] = -8'd42;
        rom[12][16] = -8'd8;
        rom[12][17] = 8'd0;
        rom[12][18] = 8'd22;
        rom[12][19] = 8'd17;
        rom[12][20] = -8'd9;
        rom[12][21] = 8'd1;
        rom[12][22] = -8'd30;
        rom[12][23] = -8'd32;
        rom[12][24] = 8'd1;
        rom[12][25] = 8'd22;
        rom[12][26] = 8'd17;
        rom[12][27] = 8'd7;
        rom[12][28] = 8'd49;
        rom[12][29] = 8'd2;
        rom[12][30] = -8'd19;
        rom[12][31] = 8'd27;
        rom[13][0] = -8'd42;
        rom[13][1] = -8'd13;
        rom[13][2] = -8'd23;
        rom[13][3] = -8'd5;
        rom[13][4] = -8'd2;
        rom[13][5] = 8'd17;
        rom[13][6] = 8'd36;
        rom[13][7] = -8'd21;
        rom[13][8] = 8'd30;
        rom[13][9] = -8'd24;
        rom[13][10] = 8'd6;
        rom[13][11] = -8'd29;
        rom[13][12] = -8'd14;
        rom[13][13] = -8'd53;
        rom[13][14] = 8'd19;
        rom[13][15] = -8'd3;
        rom[13][16] = -8'd27;
        rom[13][17] = 8'd9;
        rom[13][18] = -8'd51;
        rom[13][19] = -8'd43;
        rom[13][20] = -8'd52;
        rom[13][21] = -8'd43;
        rom[13][22] = -8'd28;
        rom[13][23] = -8'd38;
        rom[13][24] = 8'd32;
        rom[13][25] = -8'd15;
        rom[13][26] = -8'd42;
        rom[13][27] = -8'd32;
        rom[13][28] = -8'd15;
        rom[13][29] = -8'd7;
        rom[13][30] = 8'd17;
        rom[13][31] = -8'd2;
        rom[14][0] = 8'd35;
        rom[14][1] = -8'd18;
        rom[14][2] = -8'd23;
        rom[14][3] = 8'd6;
        rom[14][4] = 8'd34;
        rom[14][5] = -8'd47;
        rom[14][6] = -8'd27;
        rom[14][7] = -8'd15;
        rom[14][8] = -8'd1;
        rom[14][9] = 8'd18;
        rom[14][10] = -8'd6;
        rom[14][11] = -8'd6;
        rom[14][12] = -8'd5;
        rom[14][13] = 8'd10;
        rom[14][14] = -8'd6;
        rom[14][15] = 8'd17;
        rom[14][16] = -8'd10;
        rom[14][17] = -8'd22;
        rom[14][18] = -8'd25;
        rom[14][19] = 8'd4;
        rom[14][20] = -8'd1;
        rom[14][21] = -8'd3;
        rom[14][22] = 8'd1;
        rom[14][23] = 8'd2;
        rom[14][24] = -8'd28;
        rom[14][25] = 8'd14;
        rom[14][26] = 8'd5;
        rom[14][27] = -8'd15;
        rom[14][28] = 8'd7;
        rom[14][29] = -8'd10;
        rom[14][30] = 8'd11;
        rom[14][31] = -8'd6;
        rom[15][0] = -8'd6;
        rom[15][1] = -8'd10;
        rom[15][2] = -8'd6;
        rom[15][3] = -8'd1;
        rom[15][4] = 8'd28;
        rom[15][5] = -8'd32;
        rom[15][6] = 8'd34;
        rom[15][7] = 8'd6;
        rom[15][8] = 8'd15;
        rom[15][9] = 8'd0;
        rom[15][10] = 8'd10;
        rom[15][11] = 8'd7;
        rom[15][12] = -8'd2;
        rom[15][13] = 8'd7;
        rom[15][14] = 8'd51;
        rom[15][15] = -8'd21;
        rom[15][16] = 8'd19;
        rom[15][17] = 8'd12;
        rom[15][18] = -8'd48;
        rom[15][19] = 8'd53;
        rom[15][20] = 8'd30;
        rom[15][21] = 8'd23;
        rom[15][22] = -8'd10;
        rom[15][23] = -8'd24;
        rom[15][24] = 8'd0;
        rom[15][25] = -8'd2;
        rom[15][26] = 8'd22;
        rom[15][27] = 8'd2;
        rom[15][28] = -8'd12;
        rom[15][29] = 8'd3;
        rom[15][30] = 8'd2;
        rom[15][31] = 8'd0;
        rom[16][0] = -8'd18;
        rom[16][1] = 8'd17;
        rom[16][2] = 8'd33;
        rom[16][3] = 8'd21;
        rom[16][4] = -8'd1;
        rom[16][5] = 8'd19;
        rom[16][6] = -8'd15;
        rom[16][7] = -8'd24;
        rom[16][8] = 8'd9;
        rom[16][9] = -8'd7;
        rom[16][10] = -8'd11;
        rom[16][11] = -8'd31;
        rom[16][12] = 8'd4;
        rom[16][13] = 8'd1;
        rom[16][14] = -8'd10;
        rom[16][15] = -8'd25;
        rom[16][16] = -8'd8;
        rom[16][17] = 8'd4;
        rom[16][18] = -8'd4;
        rom[16][19] = -8'd16;
        rom[16][20] = 8'd25;
        rom[16][21] = -8'd55;
        rom[16][22] = -8'd9;
        rom[16][23] = -8'd54;
        rom[16][24] = -8'd45;
        rom[16][25] = -8'd17;
        rom[16][26] = 8'd4;
        rom[16][27] = 8'd0;
        rom[16][28] = -8'd16;
        rom[16][29] = 8'd3;
        rom[16][30] = -8'd11;
        rom[16][31] = 8'd8;
        rom[17][0] = -8'd7;
        rom[17][1] = -8'd29;
        rom[17][2] = 8'd35;
        rom[17][3] = 8'd25;
        rom[17][4] = 8'd18;
        rom[17][5] = -8'd2;
        rom[17][6] = -8'd5;
        rom[17][7] = 8'd1;
        rom[17][8] = 8'd0;
        rom[17][9] = 8'd13;
        rom[17][10] = 8'd40;
        rom[17][11] = -8'd12;
        rom[17][12] = 8'd11;
        rom[17][13] = 8'd7;
        rom[17][14] = -8'd19;
        rom[17][15] = -8'd11;
        rom[17][16] = 8'd9;
        rom[17][17] = -8'd20;
        rom[17][18] = -8'd17;
        rom[17][19] = -8'd15;
        rom[17][20] = 8'd34;
        rom[17][21] = -8'd5;
        rom[17][22] = 8'd6;
        rom[17][23] = 8'd3;
        rom[17][24] = -8'd14;
        rom[17][25] = 8'd38;
        rom[17][26] = -8'd11;
        rom[17][27] = -8'd8;
        rom[17][28] = 8'd12;
        rom[17][29] = -8'd6;
        rom[17][30] = 8'd7;
        rom[17][31] = -8'd26;
        rom[18][0] = 8'd0;
        rom[18][1] = -8'd5;
        rom[18][2] = 8'd48;
        rom[18][3] = 8'd42;
        rom[18][4] = 8'd17;
        rom[18][5] = -8'd26;
        rom[18][6] = 8'd16;
        rom[18][7] = -8'd6;
        rom[18][8] = 8'd32;
        rom[18][9] = -8'd24;
        rom[18][10] = 8'd0;
        rom[18][11] = -8'd3;
        rom[18][12] = -8'd21;
        rom[18][13] = 8'd0;
        rom[18][14] = -8'd11;
        rom[18][15] = -8'd37;
        rom[18][16] = 8'd63;
        rom[18][17] = 8'd31;
        rom[18][18] = 8'd19;
        rom[18][19] = 8'd10;
        rom[18][20] = 8'd16;
        rom[18][21] = 8'd17;
        rom[18][22] = 8'd1;
        rom[18][23] = -8'd31;
        rom[18][24] = -8'd9;
        rom[18][25] = 8'd16;
        rom[18][26] = -8'd14;
        rom[18][27] = -8'd7;
        rom[18][28] = 8'd45;
        rom[18][29] = -8'd5;
        rom[18][30] = 8'd37;
        rom[18][31] = -8'd20;
        rom[19][0] = -8'd16;
        rom[19][1] = -8'd1;
        rom[19][2] = -8'd56;
        rom[19][3] = 8'd27;
        rom[19][4] = -8'd14;
        rom[19][5] = -8'd1;
        rom[19][6] = 8'd38;
        rom[19][7] = 8'd7;
        rom[19][8] = -8'd29;
        rom[19][9] = -8'd15;
        rom[19][10] = -8'd7;
        rom[19][11] = -8'd9;
        rom[19][12] = -8'd29;
        rom[19][13] = 8'd46;
        rom[19][14] = 8'd34;
        rom[19][15] = -8'd11;
        rom[19][16] = 8'd4;
        rom[19][17] = 8'd8;
        rom[19][18] = 8'd67;
        rom[19][19] = 8'd1;
        rom[19][20] = -8'd7;
        rom[19][21] = 8'd6;
        rom[19][22] = 8'd31;
        rom[19][23] = -8'd8;
        rom[19][24] = -8'd36;
        rom[19][25] = -8'd35;
        rom[19][26] = 8'd19;
        rom[19][27] = -8'd2;
        rom[19][28] = 8'd15;
        rom[19][29] = -8'd3;
        rom[19][30] = 8'd11;
        rom[19][31] = -8'd25;
        rom[20][0] = 8'd48;
        rom[20][1] = 8'd34;
        rom[20][2] = -8'd23;
        rom[20][3] = -8'd3;
        rom[20][4] = -8'd14;
        rom[20][5] = -8'd6;
        rom[20][6] = -8'd13;
        rom[20][7] = 8'd15;
        rom[20][8] = -8'd46;
        rom[20][9] = -8'd10;
        rom[20][10] = 8'd25;
        rom[20][11] = -8'd14;
        rom[20][12] = 8'd32;
        rom[20][13] = -8'd5;
        rom[20][14] = 8'd2;
        rom[20][15] = 8'd4;
        rom[20][16] = -8'd35;
        rom[20][17] = 8'd9;
        rom[20][18] = -8'd11;
        rom[20][19] = 8'd2;
        rom[20][20] = 8'd19;
        rom[20][21] = 8'd18;
        rom[20][22] = -8'd37;
        rom[20][23] = -8'd14;
        rom[20][24] = -8'd11;
        rom[20][25] = 8'd13;
        rom[20][26] = -8'd4;
        rom[20][27] = 8'd12;
        rom[20][28] = -8'd12;
        rom[20][29] = 8'd4;
        rom[20][30] = -8'd29;
        rom[20][31] = 8'd3;
        rom[21][0] = -8'd37;
        rom[21][1] = 8'd10;
        rom[21][2] = 8'd3;
        rom[21][3] = 8'd10;
        rom[21][4] = -8'd10;
        rom[21][5] = 8'd10;
        rom[21][6] = 8'd14;
        rom[21][7] = -8'd1;
        rom[21][8] = -8'd28;
        rom[21][9] = -8'd5;
        rom[21][10] = -8'd6;
        rom[21][11] = -8'd8;
        rom[21][12] = -8'd25;
        rom[21][13] = 8'd10;
        rom[21][14] = 8'd7;
        rom[21][15] = 8'd24;
        rom[21][16] = -8'd16;
        rom[21][17] = 8'd8;
        rom[21][18] = -8'd38;
        rom[21][19] = -8'd16;
        rom[21][20] = -8'd3;
        rom[21][21] = -8'd17;
        rom[21][22] = 8'd33;
        rom[21][23] = 8'd10;
        rom[21][24] = -8'd16;
        rom[21][25] = -8'd14;
        rom[21][26] = -8'd21;
        rom[21][27] = 8'd13;
        rom[21][28] = -8'd18;
        rom[21][29] = -8'd13;
        rom[21][30] = 8'd24;
        rom[21][31] = -8'd30;
        rom[22][0] = -8'd42;
        rom[22][1] = -8'd31;
        rom[22][2] = -8'd12;
        rom[22][3] = 8'd28;
        rom[22][4] = 8'd12;
        rom[22][5] = -8'd64;
        rom[22][6] = 8'd16;
        rom[22][7] = 8'd25;
        rom[22][8] = -8'd49;
        rom[22][9] = 8'd8;
        rom[22][10] = 8'd50;
        rom[22][11] = -8'd11;
        rom[22][12] = -8'd13;
        rom[22][13] = -8'd10;
        rom[22][14] = 8'd5;
        rom[22][15] = -8'd26;
        rom[22][16] = -8'd18;
        rom[22][17] = 8'd4;
        rom[22][18] = -8'd7;
        rom[22][19] = 8'd7;
        rom[22][20] = 8'd5;
        rom[22][21] = -8'd10;
        rom[22][22] = -8'd15;
        rom[22][23] = 8'd6;
        rom[22][24] = 8'd6;
        rom[22][25] = 8'd35;
        rom[22][26] = -8'd35;
        rom[22][27] = 8'd24;
        rom[22][28] = -8'd10;
        rom[22][29] = 8'd0;
        rom[22][30] = 8'd21;
        rom[22][31] = 8'd16;
        rom[23][0] = 8'd17;
        rom[23][1] = 8'd7;
        rom[23][2] = 8'd9;
        rom[23][3] = 8'd35;
        rom[23][4] = 8'd11;
        rom[23][5] = -8'd9;
        rom[23][6] = -8'd4;
        rom[23][7] = -8'd9;
        rom[23][8] = -8'd32;
        rom[23][9] = 8'd9;
        rom[23][10] = 8'd2;
        rom[23][11] = 8'd11;
        rom[23][12] = 8'd13;
        rom[23][13] = 8'd3;
        rom[23][14] = 8'd43;
        rom[23][15] = 8'd11;
        rom[23][16] = 8'd11;
        rom[23][17] = 8'd37;
        rom[23][18] = -8'd25;
        rom[23][19] = 8'd15;
        rom[23][20] = 8'd0;
        rom[23][21] = -8'd22;
        rom[23][22] = 8'd22;
        rom[23][23] = 8'd53;
        rom[23][24] = -8'd35;
        rom[23][25] = 8'd17;
        rom[23][26] = 8'd29;
        rom[23][27] = 8'd7;
        rom[23][28] = 8'd15;
        rom[23][29] = 8'd4;
        rom[23][30] = 8'd17;
        rom[23][31] = 8'd11;
        rom[24][0] = -8'd60;
        rom[24][1] = 8'd17;
        rom[24][2] = -8'd14;
        rom[24][3] = -8'd38;
        rom[24][4] = 8'd20;
        rom[24][5] = 8'd30;
        rom[24][6] = 8'd12;
        rom[24][7] = -8'd6;
        rom[24][8] = -8'd5;
        rom[24][9] = 8'd6;
        rom[24][10] = -8'd10;
        rom[24][11] = -8'd3;
        rom[24][12] = 8'd5;
        rom[24][13] = -8'd18;
        rom[24][14] = 8'd26;
        rom[24][15] = -8'd42;
        rom[24][16] = -8'd19;
        rom[24][17] = 8'd21;
        rom[24][18] = 8'd1;
        rom[24][19] = -8'd22;
        rom[24][20] = 8'd40;
        rom[24][21] = 8'd27;
        rom[24][22] = -8'd17;
        rom[24][23] = -8'd12;
        rom[24][24] = -8'd31;
        rom[24][25] = -8'd42;
        rom[24][26] = -8'd39;
        rom[24][27] = 8'd14;
        rom[24][28] = -8'd2;
        rom[24][29] = 8'd4;
        rom[24][30] = -8'd1;
        rom[24][31] = 8'd22;
        rom[25][0] = 8'd6;
        rom[25][1] = -8'd19;
        rom[25][2] = -8'd8;
        rom[25][3] = -8'd5;
        rom[25][4] = -8'd38;
        rom[25][5] = -8'd19;
        rom[25][6] = 8'd20;
        rom[25][7] = 8'd30;
        rom[25][8] = -8'd49;
        rom[25][9] = 8'd19;
        rom[25][10] = -8'd17;
        rom[25][11] = -8'd4;
        rom[25][12] = -8'd8;
        rom[25][13] = 8'd11;
        rom[25][14] = -8'd10;
        rom[25][15] = -8'd28;
        rom[25][16] = 8'd15;
        rom[25][17] = 8'd45;
        rom[25][18] = -8'd34;
        rom[25][19] = 8'd0;
        rom[25][20] = -8'd2;
        rom[25][21] = -8'd26;
        rom[25][22] = 8'd2;
        rom[25][23] = 8'd14;
        rom[25][24] = 8'd17;
        rom[25][25] = -8'd43;
        rom[25][26] = -8'd42;
        rom[25][27] = -8'd5;
        rom[25][28] = -8'd20;
        rom[25][29] = -8'd10;
        rom[25][30] = -8'd15;
        rom[25][31] = 8'd23;
        rom[26][0] = -8'd29;
        rom[26][1] = -8'd12;
        rom[26][2] = 8'd0;
        rom[26][3] = -8'd30;
        rom[26][4] = 8'd10;
        rom[26][5] = 8'd27;
        rom[26][6] = -8'd14;
        rom[26][7] = -8'd29;
        rom[26][8] = 8'd26;
        rom[26][9] = 8'd21;
        rom[26][10] = 8'd2;
        rom[26][11] = 8'd8;
        rom[26][12] = 8'd4;
        rom[26][13] = -8'd3;
        rom[26][14] = 8'd4;
        rom[26][15] = 8'd7;
        rom[26][16] = 8'd39;
        rom[26][17] = 8'd27;
        rom[26][18] = -8'd44;
        rom[26][19] = 8'd19;
        rom[26][20] = 8'd1;
        rom[26][21] = -8'd6;
        rom[26][22] = 8'd24;
        rom[26][23] = -8'd4;
        rom[26][24] = 8'd8;
        rom[26][25] = -8'd29;
        rom[26][26] = 8'd25;
        rom[26][27] = 8'd6;
        rom[26][28] = 8'd8;
        rom[26][29] = -8'd5;
        rom[26][30] = 8'd8;
        rom[26][31] = -8'd2;
        rom[27][0] = 8'd10;
        rom[27][1] = -8'd5;
        rom[27][2] = -8'd4;
        rom[27][3] = 8'd11;
        rom[27][4] = 8'd33;
        rom[27][5] = -8'd5;
        rom[27][6] = 8'd18;
        rom[27][7] = 8'd12;
        rom[27][8] = -8'd41;
        rom[27][9] = -8'd9;
        rom[27][10] = -8'd6;
        rom[27][11] = 8'd21;
        rom[27][12] = -8'd5;
        rom[27][13] = 8'd46;
        rom[27][14] = 8'd2;
        rom[27][15] = -8'd6;
        rom[27][16] = -8'd21;
        rom[27][17] = -8'd2;
        rom[27][18] = 8'd1;
        rom[27][19] = -8'd25;
        rom[27][20] = -8'd10;
        rom[27][21] = 8'd8;
        rom[27][22] = 8'd1;
        rom[27][23] = 8'd0;
        rom[27][24] = -8'd28;
        rom[27][25] = -8'd26;
        rom[27][26] = -8'd15;
        rom[27][27] = -8'd16;
        rom[27][28] = 8'd8;
        rom[27][29] = -8'd8;
        rom[27][30] = -8'd2;
        rom[27][31] = -8'd5;
        rom[28][0] = 8'd4;
        rom[28][1] = -8'd28;
        rom[28][2] = 8'd19;
        rom[28][3] = 8'd6;
        rom[28][4] = -8'd4;
        rom[28][5] = 8'd6;
        rom[28][6] = 8'd35;
        rom[28][7] = 8'd32;
        rom[28][8] = 8'd36;
        rom[28][9] = -8'd10;
        rom[28][10] = -8'd31;
        rom[28][11] = 8'd5;
        rom[28][12] = -8'd3;
        rom[28][13] = -8'd30;
        rom[28][14] = 8'd30;
        rom[28][15] = -8'd42;
        rom[28][16] = -8'd27;
        rom[28][17] = 8'd10;
        rom[28][18] = -8'd8;
        rom[28][19] = 8'd1;
        rom[28][20] = -8'd58;
        rom[28][21] = -8'd12;
        rom[28][22] = -8'd4;
        rom[28][23] = -8'd44;
        rom[28][24] = -8'd3;
        rom[28][25] = -8'd16;
        rom[28][26] = 8'd3;
        rom[28][27] = 8'd42;
        rom[28][28] = -8'd22;
        rom[28][29] = -8'd1;
        rom[28][30] = -8'd23;
        rom[28][31] = 8'd3;
        rom[29][0] = -8'd2;
        rom[29][1] = 8'd14;
        rom[29][2] = 8'd17;
        rom[29][3] = 8'd8;
        rom[29][4] = 8'd8;
        rom[29][5] = -8'd28;
        rom[29][6] = 8'd6;
        rom[29][7] = -8'd38;
        rom[29][8] = -8'd7;
        rom[29][9] = 8'd54;
        rom[29][10] = 8'd14;
        rom[29][11] = -8'd7;
        rom[29][12] = 8'd12;
        rom[29][13] = -8'd14;
        rom[29][14] = -8'd14;
        rom[29][15] = -8'd9;
        rom[29][16] = 8'd23;
        rom[29][17] = -8'd5;
        rom[29][18] = 8'd22;
        rom[29][19] = 8'd49;
        rom[29][20] = 8'd18;
        rom[29][21] = 8'd28;
        rom[29][22] = -8'd49;
        rom[29][23] = 8'd44;
        rom[29][24] = -8'd44;
        rom[29][25] = 8'd26;
        rom[29][26] = 8'd17;
        rom[29][27] = 8'd14;
        rom[29][28] = 8'd11;
        rom[29][29] = -8'd12;
        rom[29][30] = 8'd15;
        rom[29][31] = 8'd0;
        rom[30][0] = 8'd32;
        rom[30][1] = -8'd35;
        rom[30][2] = -8'd5;
        rom[30][3] = -8'd27;
        rom[30][4] = -8'd34;
        rom[30][5] = -8'd16;
        rom[30][6] = -8'd7;
        rom[30][7] = -8'd21;
        rom[30][8] = -8'd25;
        rom[30][9] = -8'd54;
        rom[30][10] = 8'd9;
        rom[30][11] = -8'd24;
        rom[30][12] = 8'd6;
        rom[30][13] = 8'd27;
        rom[30][14] = 8'd34;
        rom[30][15] = 8'd48;
        rom[30][16] = -8'd34;
        rom[30][17] = -8'd13;
        rom[30][18] = 8'd35;
        rom[30][19] = 8'd13;
        rom[30][20] = 8'd8;
        rom[30][21] = 8'd23;
        rom[30][22] = -8'd10;
        rom[30][23] = -8'd67;
        rom[30][24] = 8'd14;
        rom[30][25] = -8'd1;
        rom[30][26] = 8'd3;
        rom[30][27] = 8'd24;
        rom[30][28] = 8'd33;
        rom[30][29] = 8'd9;
        rom[30][30] = -8'd15;
        rom[30][31] = 8'd5;
        rom[31][0] = -8'd33;
        rom[31][1] = 8'd12;
        rom[31][2] = 8'd37;
        rom[31][3] = 8'd3;
        rom[31][4] = 8'd34;
        rom[31][5] = 8'd1;
        rom[31][6] = -8'd3;
        rom[31][7] = 8'd3;
        rom[31][8] = 8'd18;
        rom[31][9] = -8'd42;
        rom[31][10] = -8'd23;
        rom[31][11] = -8'd49;
        rom[31][12] = -8'd3;
        rom[31][13] = 8'd51;
        rom[31][14] = -8'd15;
        rom[31][15] = 8'd34;
        rom[31][16] = 8'd36;
        rom[31][17] = 8'd15;
        rom[31][18] = 8'd28;
        rom[31][19] = -8'd45;
        rom[31][20] = -8'd25;
        rom[31][21] = -8'd4;
        rom[31][22] = 8'd19;
        rom[31][23] = -8'd41;
        rom[31][24] = 8'd11;
        rom[31][25] = 8'd18;
        rom[31][26] = 8'd3;
        rom[31][27] = -8'd21;
        rom[31][28] = -8'd21;
        rom[31][29] = -8'd14;
        rom[31][30] = -8'd36;
        rom[31][31] = -8'd10;
        rom[32][0] = 8'd5;
        rom[32][1] = 8'd7;
        rom[32][2] = 8'd19;
        rom[32][3] = -8'd28;
        rom[32][4] = 8'd31;
        rom[32][5] = -8'd33;
        rom[32][6] = 8'd0;
        rom[32][7] = -8'd5;
        rom[32][8] = 8'd12;
        rom[32][9] = 8'd16;
        rom[32][10] = 8'd9;
        rom[32][11] = -8'd11;
        rom[32][12] = -8'd7;
        rom[32][13] = 8'd7;
        rom[32][14] = -8'd3;
        rom[32][15] = -8'd80;
        rom[32][16] = -8'd25;
        rom[32][17] = 8'd18;
        rom[32][18] = -8'd12;
        rom[32][19] = -8'd13;
        rom[32][20] = -8'd48;
        rom[32][21] = -8'd38;
        rom[32][22] = -8'd17;
        rom[32][23] = 8'd10;
        rom[32][24] = -8'd7;
        rom[32][25] = 8'd15;
        rom[32][26] = -8'd16;
        rom[32][27] = 8'd26;
        rom[32][28] = -8'd8;
        rom[32][29] = 8'd5;
        rom[32][30] = 8'd4;
        rom[32][31] = -8'd2;
        rom[33][0] = 8'd38;
        rom[33][1] = -8'd4;
        rom[33][2] = -8'd21;
        rom[33][3] = -8'd41;
        rom[33][4] = -8'd65;
        rom[33][5] = -8'd18;
        rom[33][6] = -8'd20;
        rom[33][7] = -8'd10;
        rom[33][8] = -8'd37;
        rom[33][9] = -8'd15;
        rom[33][10] = 8'd3;
        rom[33][11] = 8'd20;
        rom[33][12] = -8'd10;
        rom[33][13] = 8'd23;
        rom[33][14] = 8'd17;
        rom[33][15] = -8'd5;
        rom[33][16] = 8'd53;
        rom[33][17] = 8'd42;
        rom[33][18] = 8'd33;
        rom[33][19] = -8'd6;
        rom[33][20] = -8'd23;
        rom[33][21] = 8'd9;
        rom[33][22] = 8'd10;
        rom[33][23] = -8'd19;
        rom[33][24] = 8'd13;
        rom[33][25] = -8'd31;
        rom[33][26] = -8'd24;
        rom[33][27] = 8'd4;
        rom[33][28] = -8'd7;
        rom[33][29] = -8'd3;
        rom[33][30] = -8'd36;
        rom[33][31] = -8'd7;
        rom[34][0] = 8'd0;
        rom[34][1] = 8'd2;
        rom[34][2] = -8'd64;
        rom[34][3] = -8'd10;
        rom[34][4] = -8'd11;
        rom[34][5] = 8'd35;
        rom[34][6] = -8'd5;
        rom[34][7] = 8'd7;
        rom[34][8] = -8'd13;
        rom[34][9] = -8'd78;
        rom[34][10] = 8'd6;
        rom[34][11] = 8'd3;
        rom[34][12] = -8'd40;
        rom[34][13] = -8'd30;
        rom[34][14] = -8'd6;
        rom[34][15] = -8'd6;
        rom[34][16] = -8'd47;
        rom[34][17] = -8'd4;
        rom[34][18] = -8'd9;
        rom[34][19] = -8'd28;
        rom[34][20] = -8'd23;
        rom[34][21] = -8'd44;
        rom[34][22] = 8'd42;
        rom[34][23] = 8'd5;
        rom[34][24] = -8'd8;
        rom[34][25] = -8'd3;
        rom[34][26] = -8'd26;
        rom[34][27] = -8'd50;
        rom[34][28] = -8'd47;
        rom[34][29] = 8'd3;
        rom[34][30] = 8'd27;
        rom[34][31] = 8'd9;
        rom[35][0] = 8'd28;
        rom[35][1] = 8'd5;
        rom[35][2] = -8'd14;
        rom[35][3] = 8'd2;
        rom[35][4] = -8'd1;
        rom[35][5] = -8'd35;
        rom[35][6] = 8'd3;
        rom[35][7] = -8'd13;
        rom[35][8] = -8'd27;
        rom[35][9] = 8'd2;
        rom[35][10] = -8'd3;
        rom[35][11] = -8'd8;
        rom[35][12] = 8'd13;
        rom[35][13] = -8'd25;
        rom[35][14] = 8'd40;
        rom[35][15] = -8'd7;
        rom[35][16] = -8'd7;
        rom[35][17] = 8'd8;
        rom[35][18] = 8'd16;
        rom[35][19] = 8'd21;
        rom[35][20] = 8'd27;
        rom[35][21] = -8'd13;
        rom[35][22] = -8'd4;
        rom[35][23] = -8'd31;
        rom[35][24] = 8'd5;
        rom[35][25] = 8'd24;
        rom[35][26] = 8'd0;
        rom[35][27] = 8'd6;
        rom[35][28] = -8'd29;
        rom[35][29] = -8'd6;
        rom[35][30] = 8'd15;
        rom[35][31] = 8'd3;
        rom[36][0] = -8'd66;
        rom[36][1] = -8'd36;
        rom[36][2] = 8'd26;
        rom[36][3] = 8'd10;
        rom[36][4] = 8'd0;
        rom[36][5] = 8'd22;
        rom[36][6] = 8'd20;
        rom[36][7] = 8'd5;
        rom[36][8] = -8'd19;
        rom[36][9] = -8'd35;
        rom[36][10] = 8'd16;
        rom[36][11] = 8'd73;
        rom[36][12] = -8'd9;
        rom[36][13] = -8'd13;
        rom[36][14] = 8'd39;
        rom[36][15] = -8'd3;
        rom[36][16] = -8'd29;
        rom[36][17] = 8'd7;
        rom[36][18] = 8'd23;
        rom[36][19] = -8'd51;
        rom[36][20] = 8'd13;
        rom[36][21] = -8'd36;
        rom[36][22] = -8'd4;
        rom[36][23] = -8'd31;
        rom[36][24] = 8'd35;
        rom[36][25] = 8'd10;
        rom[36][26] = -8'd18;
        rom[36][27] = -8'd12;
        rom[36][28] = 8'd0;
        rom[36][29] = -8'd5;
        rom[36][30] = 8'd5;
        rom[36][31] = 8'd25;
        rom[37][0] = 8'd22;
        rom[37][1] = -8'd35;
        rom[37][2] = -8'd32;
        rom[37][3] = -8'd19;
        rom[37][4] = -8'd58;
        rom[37][5] = -8'd20;
        rom[37][6] = -8'd16;
        rom[37][7] = -8'd26;
        rom[37][8] = -8'd16;
        rom[37][9] = -8'd43;
        rom[37][10] = -8'd13;
        rom[37][11] = 8'd26;
        rom[37][12] = -8'd17;
        rom[37][13] = 8'd30;
        rom[37][14] = 8'd7;
        rom[37][15] = -8'd11;
        rom[37][16] = -8'd21;
        rom[37][17] = -8'd10;
        rom[37][18] = -8'd55;
        rom[37][19] = 8'd14;
        rom[37][20] = -8'd29;
        rom[37][21] = -8'd19;
        rom[37][22] = -8'd1;
        rom[37][23] = -8'd12;
        rom[37][24] = 8'd29;
        rom[37][25] = -8'd45;
        rom[37][26] = -8'd26;
        rom[37][27] = -8'd4;
        rom[37][28] = -8'd33;
        rom[37][29] = -8'd9;
        rom[37][30] = 8'd2;
        rom[37][31] = 8'd3;
        rom[38][0] = 8'd4;
        rom[38][1] = 8'd6;
        rom[38][2] = -8'd38;
        rom[38][3] = 8'd5;
        rom[38][4] = -8'd18;
        rom[38][5] = 8'd3;
        rom[38][6] = -8'd9;
        rom[38][7] = -8'd35;
        rom[38][8] = 8'd16;
        rom[38][9] = 8'd3;
        rom[38][10] = -8'd10;
        rom[38][11] = -8'd1;
        rom[38][12] = 8'd29;
        rom[38][13] = 8'd30;
        rom[38][14] = 8'd10;
        rom[38][15] = 8'd19;
        rom[38][16] = -8'd1;
        rom[38][17] = 8'd24;
        rom[38][18] = -8'd30;
        rom[38][19] = -8'd18;
        rom[38][20] = 8'd11;
        rom[38][21] = -8'd15;
        rom[38][22] = 8'd11;
        rom[38][23] = 8'd26;
        rom[38][24] = 8'd5;
        rom[38][25] = -8'd36;
        rom[38][26] = -8'd5;
        rom[38][27] = -8'd55;
        rom[38][28] = 8'd22;
        rom[38][29] = -8'd10;
        rom[38][30] = -8'd50;
        rom[38][31] = 8'd27;
        rom[39][0] = -8'd14;
        rom[39][1] = -8'd4;
        rom[39][2] = -8'd4;
        rom[39][3] = 8'd19;
        rom[39][4] = 8'd5;
        rom[39][5] = -8'd58;
        rom[39][6] = 8'd5;
        rom[39][7] = -8'd1;
        rom[39][8] = -8'd6;
        rom[39][9] = 8'd4;
        rom[39][10] = -8'd7;
        rom[39][11] = -8'd12;
        rom[39][12] = 8'd31;
        rom[39][13] = -8'd3;
        rom[39][14] = -8'd34;
        rom[39][15] = 8'd16;
        rom[39][16] = 8'd8;
        rom[39][17] = 8'd14;
        rom[39][18] = -8'd11;
        rom[39][19] = 8'd2;
        rom[39][20] = -8'd7;
        rom[39][21] = -8'd3;
        rom[39][22] = -8'd16;
        rom[39][23] = -8'd4;
        rom[39][24] = 8'd6;
        rom[39][25] = -8'd30;
        rom[39][26] = 8'd25;
        rom[39][27] = 8'd32;
        rom[39][28] = -8'd2;
        rom[39][29] = 8'd1;
        rom[39][30] = -8'd13;
        rom[39][31] = -8'd5;
        rom[40][0] = 8'd23;
        rom[40][1] = 8'd23;
        rom[40][2] = 8'd16;
        rom[40][3] = 8'd17;
        rom[40][4] = 8'd4;
        rom[40][5] = 8'd16;
        rom[40][6] = 8'd4;
        rom[40][7] = -8'd9;
        rom[40][8] = -8'd31;
        rom[40][9] = 8'd28;
        rom[40][10] = 8'd23;
        rom[40][11] = 8'd26;
        rom[40][12] = 8'd8;
        rom[40][13] = 8'd8;
        rom[40][14] = 8'd12;
        rom[40][15] = -8'd11;
        rom[40][16] = 8'd25;
        rom[40][17] = -8'd6;
        rom[40][18] = 8'd6;
        rom[40][19] = -8'd17;
        rom[40][20] = 8'd14;
        rom[40][21] = 8'd3;
        rom[40][22] = 8'd21;
        rom[40][23] = -8'd18;
        rom[40][24] = 8'd11;
        rom[40][25] = 8'd8;
        rom[40][26] = 8'd12;
        rom[40][27] = 8'd30;
        rom[40][28] = -8'd14;
        rom[40][29] = -8'd8;
        rom[40][30] = 8'd5;
        rom[40][31] = -8'd23;
        rom[41][0] = -8'd7;
        rom[41][1] = 8'd27;
        rom[41][2] = 8'd7;
        rom[41][3] = -8'd3;
        rom[41][4] = -8'd8;
        rom[41][5] = 8'd18;
        rom[41][6] = -8'd22;
        rom[41][7] = -8'd21;
        rom[41][8] = -8'd8;
        rom[41][9] = -8'd20;
        rom[41][10] = 8'd16;
        rom[41][11] = -8'd30;
        rom[41][12] = -8'd39;
        rom[41][13] = -8'd37;
        rom[41][14] = 8'd6;
        rom[41][15] = 8'd28;
        rom[41][16] = -8'd57;
        rom[41][17] = -8'd20;
        rom[41][18] = 8'd14;
        rom[41][19] = 8'd20;
        rom[41][20] = 8'd10;
        rom[41][21] = -8'd25;
        rom[41][22] = 8'd35;
        rom[41][23] = -8'd11;
        rom[41][24] = 8'd18;
        rom[41][25] = -8'd8;
        rom[41][26] = 8'd21;
        rom[41][27] = -8'd23;
        rom[41][28] = -8'd9;
        rom[41][29] = 8'd7;
        rom[41][30] = 8'd17;
        rom[41][31] = -8'd4;
        rom[42][0] = 8'd10;
        rom[42][1] = -8'd35;
        rom[42][2] = -8'd29;
        rom[42][3] = -8'd38;
        rom[42][4] = 8'd16;
        rom[42][5] = -8'd18;
        rom[42][6] = 8'd11;
        rom[42][7] = 8'd9;
        rom[42][8] = 8'd38;
        rom[42][9] = 8'd25;
        rom[42][10] = -8'd21;
        rom[42][11] = -8'd33;
        rom[42][12] = -8'd7;
        rom[42][13] = -8'd12;
        rom[42][14] = 8'd32;
        rom[42][15] = 8'd16;
        rom[42][16] = 8'd20;
        rom[42][17] = 8'd48;
        rom[42][18] = -8'd26;
        rom[42][19] = 8'd4;
        rom[42][20] = 8'd4;
        rom[42][21] = 8'd16;
        rom[42][22] = 8'd31;
        rom[42][23] = 8'd9;
        rom[42][24] = 8'd38;
        rom[42][25] = -8'd81;
        rom[42][26] = 8'd14;
        rom[42][27] = -8'd43;
        rom[42][28] = -8'd5;
        rom[42][29] = 8'd0;
        rom[42][30] = 8'd34;
        rom[42][31] = -8'd7;
        rom[43][0] = -8'd14;
        rom[43][1] = 8'd0;
        rom[43][2] = -8'd35;
        rom[43][3] = -8'd20;
        rom[43][4] = -8'd13;
        rom[43][5] = -8'd26;
        rom[43][6] = 8'd7;
        rom[43][7] = 8'd13;
        rom[43][8] = -8'd24;
        rom[43][9] = -8'd20;
        rom[43][10] = 8'd0;
        rom[43][11] = -8'd15;
        rom[43][12] = 8'd26;
        rom[43][13] = -8'd4;
        rom[43][14] = 8'd23;
        rom[43][15] = 8'd17;
        rom[43][16] = -8'd5;
        rom[43][17] = 8'd14;
        rom[43][18] = 8'd31;
        rom[43][19] = 8'd25;
        rom[43][20] = 8'd16;
        rom[43][21] = 8'd32;
        rom[43][22] = -8'd13;
        rom[43][23] = 8'd31;
        rom[43][24] = 8'd27;
        rom[43][25] = -8'd41;
        rom[43][26] = 8'd3;
        rom[43][27] = -8'd10;
        rom[43][28] = 8'd4;
        rom[43][29] = -8'd13;
        rom[43][30] = -8'd11;
        rom[43][31] = -8'd4;
        rom[44][0] = 8'd58;
        rom[44][1] = 8'd4;
        rom[44][2] = 8'd1;
        rom[44][3] = -8'd8;
        rom[44][4] = -8'd22;
        rom[44][5] = -8'd3;
        rom[44][6] = -8'd1;
        rom[44][7] = -8'd28;
        rom[44][8] = -8'd4;
        rom[44][9] = -8'd27;
        rom[44][10] = 8'd25;
        rom[44][11] = -8'd17;
        rom[44][12] = -8'd4;
        rom[44][13] = -8'd12;
        rom[44][14] = 8'd23;
        rom[44][15] = -8'd28;
        rom[44][16] = 8'd20;
        rom[44][17] = -8'd2;
        rom[44][18] = 8'd8;
        rom[44][19] = 8'd2;
        rom[44][20] = -8'd1;
        rom[44][21] = -8'd23;
        rom[44][22] = -8'd23;
        rom[44][23] = -8'd10;
        rom[44][24] = 8'd19;
        rom[44][25] = 8'd38;
        rom[44][26] = 8'd20;
        rom[44][27] = 8'd3;
        rom[44][28] = -8'd8;
        rom[44][29] = -8'd1;
        rom[44][30] = -8'd52;
        rom[44][31] = 8'd3;
        rom[45][0] = 8'd4;
        rom[45][1] = -8'd33;
        rom[45][2] = -8'd24;
        rom[45][3] = -8'd37;
        rom[45][4] = -8'd16;
        rom[45][5] = 8'd61;
        rom[45][6] = 8'd8;
        rom[45][7] = -8'd17;
        rom[45][8] = -8'd34;
        rom[45][9] = -8'd54;
        rom[45][10] = 8'd43;
        rom[45][11] = -8'd21;
        rom[45][12] = 8'd6;
        rom[45][13] = -8'd58;
        rom[45][14] = 8'd11;
        rom[45][15] = 8'd7;
        rom[45][16] = -8'd20;
        rom[45][17] = -8'd5;
        rom[45][18] = -8'd43;
        rom[45][19] = -8'd16;
        rom[45][20] = -8'd42;
        rom[45][21] = -8'd58;
        rom[45][22] = -8'd22;
        rom[45][23] = -8'd7;
        rom[45][24] = 8'd32;
        rom[45][25] = 8'd9;
        rom[45][26] = -8'd46;
        rom[45][27] = -8'd36;
        rom[45][28] = -8'd31;
        rom[45][29] = -8'd6;
        rom[45][30] = -8'd6;
        rom[45][31] = -8'd3;
        rom[46][0] = 8'd12;
        rom[46][1] = 8'd9;
        rom[46][2] = 8'd19;
        rom[46][3] = 8'd18;
        rom[46][4] = 8'd24;
        rom[46][5] = -8'd56;
        rom[46][6] = -8'd9;
        rom[46][7] = -8'd6;
        rom[46][8] = 8'd1;
        rom[46][9] = 8'd15;
        rom[46][10] = 8'd14;
        rom[46][11] = 8'd10;
        rom[46][12] = -8'd14;
        rom[46][13] = -8'd19;
        rom[46][14] = -8'd18;
        rom[46][15] = 8'd7;
        rom[46][16] = -8'd26;
        rom[46][17] = -8'd12;
        rom[46][18] = 8'd0;
        rom[46][19] = -8'd1;
        rom[46][20] = 8'd7;
        rom[46][21] = -8'd20;
        rom[46][22] = -8'd28;
        rom[46][23] = -8'd7;
        rom[46][24] = -8'd22;
        rom[46][25] = 8'd23;
        rom[46][26] = -8'd3;
        rom[46][27] = -8'd7;
        rom[46][28] = 8'd9;
        rom[46][29] = -8'd10;
        rom[46][30] = -8'd9;
        rom[46][31] = -8'd18;
        rom[47][0] = 8'd6;
        rom[47][1] = 8'd22;
        rom[47][2] = -8'd17;
        rom[47][3] = 8'd2;
        rom[47][4] = 8'd19;
        rom[47][5] = 8'd27;
        rom[47][6] = 8'd27;
        rom[47][7] = 8'd1;
        rom[47][8] = -8'd7;
        rom[47][9] = -8'd25;
        rom[47][10] = -8'd22;
        rom[47][11] = 8'd15;
        rom[47][12] = -8'd30;
        rom[47][13] = -8'd30;
        rom[47][14] = -8'd44;
        rom[47][15] = -8'd3;
        rom[47][16] = 8'd12;
        rom[47][17] = 8'd8;
        rom[47][18] = -8'd47;
        rom[47][19] = 8'd41;
        rom[47][20] = -8'd10;
        rom[47][21] = -8'd18;
        rom[47][22] = -8'd12;
        rom[47][23] = -8'd7;
        rom[47][24] = 8'd13;
        rom[47][25] = -8'd7;
        rom[47][26] = 8'd17;
        rom[47][27] = 8'd9;
        rom[47][28] = -8'd10;
        rom[47][29] = 8'd0;
        rom[47][30] = 8'd4;
        rom[47][31] = 8'd35;
        rom[48][0] = -8'd9;
        rom[48][1] = 8'd13;
        rom[48][2] = 8'd24;
        rom[48][3] = 8'd21;
        rom[48][4] = -8'd14;
        rom[48][5] = 8'd37;
        rom[48][6] = -8'd23;
        rom[48][7] = 8'd10;
        rom[48][8] = 8'd2;
        rom[48][9] = 8'd15;
        rom[48][10] = -8'd6;
        rom[48][11] = 8'd5;
        rom[48][12] = 8'd28;
        rom[48][13] = 8'd8;
        rom[48][14] = 8'd11;
        rom[48][15] = -8'd21;
        rom[48][16] = -8'd4;
        rom[48][17] = -8'd25;
        rom[48][18] = 8'd11;
        rom[48][19] = -8'd48;
        rom[48][20] = 8'd23;
        rom[48][21] = -8'd48;
        rom[48][22] = 8'd9;
        rom[48][23] = -8'd14;
        rom[48][24] = 8'd11;
        rom[48][25] = -8'd15;
        rom[48][26] = 8'd6;
        rom[48][27] = -8'd14;
        rom[48][28] = -8'd20;
        rom[48][29] = 8'd6;
        rom[48][30] = -8'd16;
        rom[48][31] = -8'd21;
        rom[49][0] = -8'd29;
        rom[49][1] = -8'd27;
        rom[49][2] = 8'd17;
        rom[49][3] = 8'd25;
        rom[49][4] = -8'd6;
        rom[49][5] = -8'd37;
        rom[49][6] = 8'd11;
        rom[49][7] = 8'd37;
        rom[49][8] = -8'd17;
        rom[49][9] = 8'd10;
        rom[49][10] = 8'd26;
        rom[49][11] = 8'd2;
        rom[49][12] = -8'd24;
        rom[49][13] = -8'd15;
        rom[49][14] = -8'd25;
        rom[49][15] = -8'd22;
        rom[49][16] = -8'd59;
        rom[49][17] = -8'd4;
        rom[49][18] = -8'd37;
        rom[49][19] = 8'd4;
        rom[49][20] = -8'd17;
        rom[49][21] = -8'd34;
        rom[49][22] = -8'd7;
        rom[49][23] = 8'd27;
        rom[49][24] = 8'd8;
        rom[49][25] = 8'd12;
        rom[49][26] = 8'd14;
        rom[49][27] = -8'd19;
        rom[49][28] = 8'd9;
        rom[49][29] = -8'd10;
        rom[49][30] = -8'd2;
        rom[49][31] = -8'd1;
        rom[50][0] = 8'd24;
        rom[50][1] = -8'd15;
        rom[50][2] = 8'd50;
        rom[50][3] = 8'd22;
        rom[50][4] = 8'd41;
        rom[50][5] = 8'd19;
        rom[50][6] = 8'd9;
        rom[50][7] = 8'd4;
        rom[50][8] = 8'd27;
        rom[50][9] = -8'd27;
        rom[50][10] = 8'd15;
        rom[50][11] = 8'd6;
        rom[50][12] = -8'd5;
        rom[50][13] = -8'd41;
        rom[50][14] = -8'd33;
        rom[50][15] = -8'd83;
        rom[50][16] = -8'd35;
        rom[50][17] = -8'd4;
        rom[50][18] = -8'd46;
        rom[50][19] = -8'd29;
        rom[50][20] = 8'd22;
        rom[50][21] = -8'd23;
        rom[50][22] = 8'd12;
        rom[50][23] = -8'd34;
        rom[50][24] = 8'd0;
        rom[50][25] = 8'd51;
        rom[50][26] = -8'd3;
        rom[50][27] = -8'd16;
        rom[50][28] = 8'd41;
        rom[50][29] = 8'd2;
        rom[50][30] = 8'd29;
        rom[50][31] = 8'd10;
        rom[51][0] = 8'd25;
        rom[51][1] = -8'd35;
        rom[51][2] = -8'd3;
        rom[51][3] = 8'd23;
        rom[51][4] = -8'd16;
        rom[51][5] = -8'd2;
        rom[51][6] = 8'd22;
        rom[51][7] = 8'd3;
        rom[51][8] = -8'd24;
        rom[51][9] = -8'd33;
        rom[51][10] = 8'd5;
        rom[51][11] = -8'd3;
        rom[51][12] = -8'd44;
        rom[51][13] = 8'd14;
        rom[51][14] = 8'd16;
        rom[51][15] = 8'd14;
        rom[51][16] = 8'd7;
        rom[51][17] = 8'd3;
        rom[51][18] = 8'd50;
        rom[51][19] = 8'd7;
        rom[51][20] = 8'd11;
        rom[51][21] = -8'd2;
        rom[51][22] = 8'd19;
        rom[51][23] = -8'd58;
        rom[51][24] = -8'd30;
        rom[51][25] = -8'd24;
        rom[51][26] = -8'd24;
        rom[51][27] = 8'd11;
        rom[51][28] = -8'd1;
        rom[51][29] = -8'd8;
        rom[51][30] = 8'd18;
        rom[51][31] = -8'd25;
        rom[52][0] = -8'd3;
        rom[52][1] = 8'd5;
        rom[52][2] = -8'd21;
        rom[52][3] = -8'd14;
        rom[52][4] = -8'd29;
        rom[52][5] = 8'd10;
        rom[52][6] = 8'd3;
        rom[52][7] = 8'd14;
        rom[52][8] = -8'd32;
        rom[52][9] = 8'd4;
        rom[52][10] = -8'd4;
        rom[52][11] = -8'd34;
        rom[52][12] = 8'd15;
        rom[52][13] = 8'd6;
        rom[52][14] = -8'd24;
        rom[52][15] = 8'd20;
        rom[52][16] = -8'd38;
        rom[52][17] = 8'd20;
        rom[52][18] = -8'd19;
        rom[52][19] = -8'd11;
        rom[52][20] = 8'd21;
        rom[52][21] = 8'd31;
        rom[52][22] = -8'd32;
        rom[52][23] = 8'd15;
        rom[52][24] = -8'd15;
        rom[52][25] = -8'd2;
        rom[52][26] = 8'd29;
        rom[52][27] = 8'd11;
        rom[52][28] = -8'd12;
        rom[52][29] = -8'd10;
        rom[52][30] = -8'd30;
        rom[52][31] = -8'd13;
        rom[53][0] = -8'd77;
        rom[53][1] = -8'd35;
        rom[53][2] = -8'd47;
        rom[53][3] = -8'd16;
        rom[53][4] = 8'd7;
        rom[53][5] = -8'd39;
        rom[53][6] = 8'd24;
        rom[53][7] = 8'd4;
        rom[53][8] = -8'd18;
        rom[53][9] = -8'd28;
        rom[53][10] = -8'd6;
        rom[53][11] = 8'd0;
        rom[53][12] = -8'd10;
        rom[53][13] = 8'd8;
        rom[53][14] = 8'd5;
        rom[53][15] = 8'd21;
        rom[53][16] = -8'd11;
        rom[53][17] = -8'd1;
        rom[53][18] = 8'd2;
        rom[53][19] = 8'd20;
        rom[53][20] = -8'd7;
        rom[53][21] = -8'd15;
        rom[53][22] = 8'd28;
        rom[53][23] = -8'd2;
        rom[53][24] = 8'd12;
        rom[53][25] = -8'd56;
        rom[53][26] = -8'd12;
        rom[53][27] = 8'd3;
        rom[53][28] = -8'd35;
        rom[53][29] = -8'd7;
        rom[53][30] = -8'd47;
        rom[53][31] = -8'd41;
        rom[54][0] = -8'd60;
        rom[54][1] = 8'd8;
        rom[54][2] = 8'd4;
        rom[54][3] = 8'd38;
        rom[54][4] = -8'd18;
        rom[54][5] = -8'd74;
        rom[54][6] = -8'd4;
        rom[54][7] = 8'd28;
        rom[54][8] = -8'd4;
        rom[54][9] = 8'd30;
        rom[54][10] = 8'd42;
        rom[54][11] = 8'd5;
        rom[54][12] = 8'd7;
        rom[54][13] = -8'd10;
        rom[54][14] = 8'd7;
        rom[54][15] = -8'd10;
        rom[54][16] = 8'd11;
        rom[54][17] = 8'd32;
        rom[54][18] = -8'd7;
        rom[54][19] = 8'd7;
        rom[54][20] = 8'd4;
        rom[54][21] = -8'd21;
        rom[54][22] = -8'd13;
        rom[54][23] = 8'd9;
        rom[54][24] = 8'd16;
        rom[54][25] = 8'd7;
        rom[54][26] = -8'd9;
        rom[54][27] = 8'd8;
        rom[54][28] = 8'd6;
        rom[54][29] = -8'd1;
        rom[54][30] = 8'd9;
        rom[54][31] = 8'd13;
        rom[55][0] = 8'd8;
        rom[55][1] = 8'd10;
        rom[55][2] = 8'd6;
        rom[55][3] = 8'd17;
        rom[55][4] = 8'd8;
        rom[55][5] = 8'd17;
        rom[55][6] = -8'd3;
        rom[55][7] = 8'd7;
        rom[55][8] = -8'd27;
        rom[55][9] = 8'd4;
        rom[55][10] = -8'd18;
        rom[55][11] = 8'd15;
        rom[55][12] = -8'd22;
        rom[55][13] = 8'd8;
        rom[55][14] = 8'd3;
        rom[55][15] = 8'd29;
        rom[55][16] = -8'd9;
        rom[55][17] = 8'd36;
        rom[55][18] = -8'd13;
        rom[55][19] = 8'd2;
        rom[55][20] = 8'd7;
        rom[55][21] = 8'd0;
        rom[55][22] = 8'd28;
        rom[55][23] = 8'd13;
        rom[55][24] = -8'd43;
        rom[55][25] = -8'd85;
        rom[55][26] = 8'd17;
        rom[55][27] = 8'd27;
        rom[55][28] = 8'd23;
        rom[55][29] = -8'd6;
        rom[55][30] = 8'd6;
        rom[55][31] = 8'd1;
        rom[56][0] = 8'd12;
        rom[56][1] = -8'd25;
        rom[56][2] = -8'd31;
        rom[56][3] = -8'd42;
        rom[56][4] = 8'd36;
        rom[56][5] = 8'd51;
        rom[56][6] = -8'd1;
        rom[56][7] = -8'd13;
        rom[56][8] = -8'd5;
        rom[56][9] = -8'd24;
        rom[56][10] = 8'd31;
        rom[56][11] = 8'd40;
        rom[56][12] = 8'd46;
        rom[56][13] = 8'd20;
        rom[56][14] = 8'd27;
        rom[56][15] = -8'd23;
        rom[56][16] = -8'd17;
        rom[56][17] = -8'd72;
        rom[56][18] = 8'd3;
        rom[56][19] = -8'd21;
        rom[56][20] = -8'd2;
        rom[56][21] = -8'd26;
        rom[56][22] = -8'd21;
        rom[56][23] = -8'd35;
        rom[56][24] = -8'd2;
        rom[56][25] = -8'd46;
        rom[56][26] = -8'd50;
        rom[56][27] = -8'd23;
        rom[56][28] = -8'd9;
        rom[56][29] = 8'd3;
        rom[56][30] = -8'd16;
        rom[56][31] = 8'd12;
        rom[57][0] = 8'd24;
        rom[57][1] = -8'd8;
        rom[57][2] = -8'd22;
        rom[57][3] = -8'd5;
        rom[57][4] = -8'd18;
        rom[57][5] = -8'd30;
        rom[57][6] = 8'd1;
        rom[57][7] = 8'd15;
        rom[57][8] = -8'd21;
        rom[57][9] = 8'd19;
        rom[57][10] = -8'd35;
        rom[57][11] = -8'd1;
        rom[57][12] = -8'd7;
        rom[57][13] = 8'd47;
        rom[57][14] = 8'd6;
        rom[57][15] = -8'd17;
        rom[57][16] = 8'd2;
        rom[57][17] = 8'd8;
        rom[57][18] = -8'd12;
        rom[57][19] = 8'd7;
        rom[57][20] = -8'd11;
        rom[57][21] = -8'd7;
        rom[57][22] = 8'd2;
        rom[57][23] = -8'd27;
        rom[57][24] = 8'd36;
        rom[57][25] = -8'd47;
        rom[57][26] = -8'd17;
        rom[57][27] = -8'd10;
        rom[57][28] = 8'd15;
        rom[57][29] = 8'd3;
        rom[57][30] = 8'd3;
        rom[57][31] = 8'd12;
        rom[58][0] = -8'd22;
        rom[58][1] = -8'd24;
        rom[58][2] = -8'd16;
        rom[58][3] = -8'd44;
        rom[58][4] = 8'd16;
        rom[58][5] = 8'd36;
        rom[58][6] = -8'd30;
        rom[58][7] = -8'd33;
        rom[58][8] = 8'd5;
        rom[58][9] = 8'd16;
        rom[58][10] = -8'd27;
        rom[58][11] = 8'd21;
        rom[58][12] = 8'd8;
        rom[58][13] = -8'd8;
        rom[58][14] = -8'd26;
        rom[58][15] = -8'd4;
        rom[58][16] = 8'd3;
        rom[58][17] = -8'd15;
        rom[58][18] = -8'd66;
        rom[58][19] = 8'd22;
        rom[58][20] = 8'd9;
        rom[58][21] = 8'd22;
        rom[58][22] = 8'd12;
        rom[58][23] = -8'd2;
        rom[58][24] = -8'd1;
        rom[58][25] = -8'd33;
        rom[58][26] = 8'd34;
        rom[58][27] = -8'd24;
        rom[58][28] = 8'd6;
        rom[58][29] = 8'd6;
        rom[58][30] = -8'd22;
        rom[58][31] = -8'd7;
        rom[59][0] = 8'd11;
        rom[59][1] = 8'd5;
        rom[59][2] = -8'd8;
        rom[59][3] = 8'd5;
        rom[59][4] = 8'd35;
        rom[59][5] = -8'd44;
        rom[59][6] = 8'd22;
        rom[59][7] = -8'd1;
        rom[59][8] = -8'd17;
        rom[59][9] = -8'd9;
        rom[59][10] = -8'd5;
        rom[59][11] = 8'd13;
        rom[59][12] = 8'd25;
        rom[59][13] = 8'd12;
        rom[59][14] = -8'd15;
        rom[59][15] = 8'd10;
        rom[59][16] = -8'd13;
        rom[59][17] = -8'd16;
        rom[59][18] = 8'd20;
        rom[59][19] = -8'd18;
        rom[59][20] = -8'd23;
        rom[59][21] = -8'd7;
        rom[59][22] = -8'd7;
        rom[59][23] = -8'd9;
        rom[59][24] = -8'd7;
        rom[59][25] = -8'd14;
        rom[59][26] = -8'd9;
        rom[59][27] = 8'd2;
        rom[59][28] = -8'd9;
        rom[59][29] = -8'd13;
        rom[59][30] = 8'd5;
        rom[59][31] = 8'd1;
        rom[60][0] = -8'd4;
        rom[60][1] = -8'd2;
        rom[60][2] = 8'd38;
        rom[60][3] = 8'd27;
        rom[60][4] = 8'd2;
        rom[60][5] = -8'd9;
        rom[60][6] = -8'd9;
        rom[60][7] = 8'd24;
        rom[60][8] = 8'd4;
        rom[60][9] = -8'd13;
        rom[60][10] = 8'd3;
        rom[60][11] = 8'd5;
        rom[60][12] = 8'd19;
        rom[60][13] = -8'd44;
        rom[60][14] = 8'd13;
        rom[60][15] = -8'd35;
        rom[60][16] = 8'd5;
        rom[60][17] = 8'd15;
        rom[60][18] = 8'd3;
        rom[60][19] = 8'd18;
        rom[60][20] = -8'd14;
        rom[60][21] = -8'd4;
        rom[60][22] = 8'd8;
        rom[60][23] = -8'd3;
        rom[60][24] = 8'd17;
        rom[60][25] = -8'd3;
        rom[60][26] = 8'd27;
        rom[60][27] = -8'd4;
        rom[60][28] = 8'd2;
        rom[60][29] = -8'd2;
        rom[60][30] = 8'd17;
        rom[60][31] = -8'd1;
        rom[61][0] = -8'd35;
        rom[61][1] = -8'd32;
        rom[61][2] = -8'd6;
        rom[61][3] = -8'd13;
        rom[61][4] = 8'd13;
        rom[61][5] = 8'd7;
        rom[61][6] = 8'd24;
        rom[61][7] = -8'd30;
        rom[61][8] = -8'd7;
        rom[61][9] = 8'd44;
        rom[61][10] = 8'd12;
        rom[61][11] = -8'd21;
        rom[61][12] = -8'd15;
        rom[61][13] = 8'd24;
        rom[61][14] = 8'd10;
        rom[61][15] = 8'd1;
        rom[61][16] = 8'd27;
        rom[61][17] = 8'd0;
        rom[61][18] = 8'd5;
        rom[61][19] = 8'd36;
        rom[61][20] = 8'd27;
        rom[61][21] = 8'd29;
        rom[61][22] = -8'd54;
        rom[61][23] = 8'd3;
        rom[61][24] = -8'd51;
        rom[61][25] = 8'd12;
        rom[61][26] = -8'd6;
        rom[61][27] = 8'd8;
        rom[61][28] = 8'd14;
        rom[61][29] = 8'd1;
        rom[61][30] = 8'd6;
        rom[61][31] = -8'd22;
        rom[62][0] = -8'd52;
        rom[62][1] = 8'd47;
        rom[62][2] = 8'd21;
        rom[62][3] = -8'd22;
        rom[62][4] = -8'd46;
        rom[62][5] = 8'd16;
        rom[62][6] = -8'd34;
        rom[62][7] = -8'd32;
        rom[62][8] = -8'd17;
        rom[62][9] = -8'd67;
        rom[62][10] = -8'd21;
        rom[62][11] = -8'd21;
        rom[62][12] = 8'd6;
        rom[62][13] = -8'd19;
        rom[62][14] = 8'd9;
        rom[62][15] = 8'd37;
        rom[62][16] = 8'd11;
        rom[62][17] = -8'd40;
        rom[62][18] = -8'd32;
        rom[62][19] = -8'd7;
        rom[62][20] = 8'd11;
        rom[62][21] = 8'd24;
        rom[62][22] = -8'd17;
        rom[62][23] = -8'd31;
        rom[62][24] = 8'd0;
        rom[62][25] = 8'd45;
        rom[62][26] = 8'd13;
        rom[62][27] = 8'd10;
        rom[62][28] = -8'd15;
        rom[62][29] = 8'd4;
        rom[62][30] = -8'd20;
        rom[62][31] = 8'd6;
        rom[63][0] = -8'd12;
        rom[63][1] = -8'd2;
        rom[63][2] = 8'd8;
        rom[63][3] = 8'd21;
        rom[63][4] = 8'd16;
        rom[63][5] = -8'd6;
        rom[63][6] = 8'd9;
        rom[63][7] = 8'd5;
        rom[63][8] = 8'd9;
        rom[63][9] = -8'd59;
        rom[63][10] = -8'd17;
        rom[63][11] = -8'd23;
        rom[63][12] = -8'd50;
        rom[63][13] = -8'd10;
        rom[63][14] = -8'd53;
        rom[63][15] = 8'd7;
        rom[63][16] = -8'd16;
        rom[63][17] = 8'd11;
        rom[63][18] = 8'd28;
        rom[63][19] = -8'd9;
        rom[63][20] = -8'd30;
        rom[63][21] = -8'd28;
        rom[63][22] = 8'd75;
        rom[63][23] = -8'd29;
        rom[63][24] = 8'd9;
        rom[63][25] = -8'd5;
        rom[63][26] = -8'd11;
        rom[63][27] = -8'd61;
        rom[63][28] = -8'd39;
        rom[63][29] = 8'd0;
        rom[63][30] = 8'd21;
        rom[63][31] = -8'd19;
        rom[64][0] = 8'd1;
        rom[64][1] = -8'd4;
        rom[64][2] = -8'd27;
        rom[64][3] = -8'd27;
        rom[64][4] = 8'd40;
        rom[64][5] = -8'd40;
        rom[64][6] = 8'd14;
        rom[64][7] = -8'd31;
        rom[64][8] = -8'd7;
        rom[64][9] = 8'd29;
        rom[64][10] = -8'd12;
        rom[64][11] = -8'd11;
        rom[64][12] = 8'd11;
        rom[64][13] = 8'd32;
        rom[64][14] = 8'd6;
        rom[64][15] = -8'd16;
        rom[64][16] = -8'd63;
        rom[64][17] = 8'd2;
        rom[64][18] = 8'd19;
        rom[64][19] = -8'd11;
        rom[64][20] = -8'd47;
        rom[64][21] = -8'd20;
        rom[64][22] = -8'd6;
        rom[64][23] = 8'd38;
        rom[64][24] = -8'd9;
        rom[64][25] = 8'd1;
        rom[64][26] = -8'd14;
        rom[64][27] = 8'd17;
        rom[64][28] = -8'd4;
        rom[64][29] = 8'd2;
        rom[64][30] = -8'd10;
        rom[64][31] = 8'd33;
        rom[65][0] = 8'd12;
        rom[65][1] = -8'd13;
        rom[65][2] = 8'd0;
        rom[65][3] = -8'd77;
        rom[65][4] = -8'd34;
        rom[65][5] = -8'd50;
        rom[65][6] = 8'd15;
        rom[65][7] = 8'd17;
        rom[65][8] = 8'd1;
        rom[65][9] = -8'd14;
        rom[65][10] = 8'd5;
        rom[65][11] = 8'd15;
        rom[65][12] = 8'd12;
        rom[65][13] = -8'd22;
        rom[65][14] = 8'd29;
        rom[65][15] = 8'd13;
        rom[65][16] = 8'd38;
        rom[65][17] = 8'd19;
        rom[65][18] = 8'd39;
        rom[65][19] = -8'd2;
        rom[65][20] = -8'd29;
        rom[65][21] = 8'd25;
        rom[65][22] = 8'd13;
        rom[65][23] = -8'd36;
        rom[65][24] = 8'd45;
        rom[65][25] = -8'd17;
        rom[65][26] = 8'd1;
        rom[65][27] = 8'd14;
        rom[65][28] = 8'd1;
        rom[65][29] = 8'd1;
        rom[65][30] = 8'd13;
        rom[65][31] = -8'd24;
        rom[66][0] = 8'd27;
        rom[66][1] = -8'd44;
        rom[66][2] = -8'd92;
        rom[66][3] = -8'd2;
        rom[66][4] = 8'd1;
        rom[66][5] = 8'd0;
        rom[66][6] = 8'd22;
        rom[66][7] = -8'd73;
        rom[66][8] = -8'd58;
        rom[66][9] = -8'd20;
        rom[66][10] = 8'd20;
        rom[66][11] = 8'd15;
        rom[66][12] = -8'd34;
        rom[66][13] = 8'd21;
        rom[66][14] = -8'd38;
        rom[66][15] = 8'd8;
        rom[66][16] = -8'd2;
        rom[66][17] = 8'd31;
        rom[66][18] = 8'd23;
        rom[66][19] = -8'd37;
        rom[66][20] = -8'd16;
        rom[66][21] = -8'd4;
        rom[66][22] = 8'd13;
        rom[66][23] = 8'd39;
        rom[66][24] = 8'd13;
        rom[66][25] = -8'd65;
        rom[66][26] = -8'd33;
        rom[66][27] = 8'd13;
        rom[66][28] = -8'd49;
        rom[66][29] = 8'd3;
        rom[66][30] = -8'd8;
        rom[66][31] = 8'd10;
        rom[67][0] = 8'd16;
        rom[67][1] = 8'd21;
        rom[67][2] = -8'd33;
        rom[67][3] = 8'd10;
        rom[67][4] = 8'd2;
        rom[67][5] = -8'd8;
        rom[67][6] = -8'd6;
        rom[67][7] = -8'd15;
        rom[67][8] = -8'd26;
        rom[67][9] = 8'd7;
        rom[67][10] = -8'd21;
        rom[67][11] = -8'd31;
        rom[67][12] = 8'd29;
        rom[67][13] = -8'd13;
        rom[67][14] = 8'd34;
        rom[67][15] = 8'd33;
        rom[67][16] = 8'd17;
        rom[67][17] = 8'd15;
        rom[67][18] = 8'd12;
        rom[67][19] = 8'd16;
        rom[67][20] = 8'd32;
        rom[67][21] = 8'd13;
        rom[67][22] = 8'd1;
        rom[67][23] = 8'd6;
        rom[67][24] = -8'd5;
        rom[67][25] = 8'd20;
        rom[67][26] = -8'd3;
        rom[67][27] = -8'd12;
        rom[67][28] = 8'd1;
        rom[67][29] = 8'd2;
        rom[67][30] = 8'd8;
        rom[67][31] = -8'd7;
        rom[68][0] = -8'd46;
        rom[68][1] = 8'd25;
        rom[68][2] = -8'd5;
        rom[68][3] = 8'd23;
        rom[68][4] = -8'd12;
        rom[68][5] = 8'd2;
        rom[68][6] = -8'd11;
        rom[68][7] = 8'd71;
        rom[68][8] = -8'd15;
        rom[68][9] = -8'd8;
        rom[68][10] = -8'd2;
        rom[68][11] = 8'd34;
        rom[68][12] = 8'd28;
        rom[68][13] = -8'd51;
        rom[68][14] = 8'd38;
        rom[68][15] = 8'd50;
        rom[68][16] = -8'd6;
        rom[68][17] = -8'd44;
        rom[68][18] = 8'd10;
        rom[68][19] = -8'd6;
        rom[68][20] = 8'd20;
        rom[68][21] = 8'd16;
        rom[68][22] = -8'd33;
        rom[68][23] = 8'd8;
        rom[68][24] = 8'd45;
        rom[68][25] = 8'd12;
        rom[68][26] = 8'd11;
        rom[68][27] = -8'd30;
        rom[68][28] = -8'd11;
        rom[68][29] = -8'd12;
        rom[68][30] = 8'd22;
        rom[68][31] = 8'd19;
        rom[69][0] = 8'd85;
        rom[69][1] = -8'd43;
        rom[69][2] = 8'd1;
        rom[69][3] = -8'd24;
        rom[69][4] = -8'd59;
        rom[69][5] = 8'd2;
        rom[69][6] = 8'd18;
        rom[69][7] = -8'd65;
        rom[69][8] = -8'd27;
        rom[69][9] = -8'd7;
        rom[69][10] = -8'd17;
        rom[69][11] = 8'd31;
        rom[69][12] = -8'd3;
        rom[69][13] = 8'd20;
        rom[69][14] = 8'd24;
        rom[69][15] = 8'd40;
        rom[69][16] = 8'd13;
        rom[69][17] = 8'd5;
        rom[69][18] = 8'd3;
        rom[69][19] = 8'd4;
        rom[69][20] = 8'd8;
        rom[69][21] = 8'd25;
        rom[69][22] = -8'd1;
        rom[69][23] = 8'd13;
        rom[69][24] = -8'd27;
        rom[69][25] = -8'd68;
        rom[69][26] = -8'd15;
        rom[69][27] = 8'd28;
        rom[69][28] = -8'd58;
        rom[69][29] = -8'd2;
        rom[69][30] = 8'd2;
        rom[69][31] = 8'd17;
        rom[70][0] = 8'd27;
        rom[70][1] = 8'd10;
        rom[70][2] = -8'd14;
        rom[70][3] = 8'd1;
        rom[70][4] = 8'd7;
        rom[70][5] = -8'd48;
        rom[70][6] = -8'd22;
        rom[70][7] = -8'd29;
        rom[70][8] = -8'd20;
        rom[70][9] = 8'd5;
        rom[70][10] = -8'd13;
        rom[70][11] = -8'd22;
        rom[70][12] = 8'd31;
        rom[70][13] = 8'd57;
        rom[70][14] = -8'd12;
        rom[70][15] = 8'd11;
        rom[70][16] = -8'd14;
        rom[70][17] = 8'd21;
        rom[70][18] = -8'd11;
        rom[70][19] = 8'd3;
        rom[70][20] = 8'd7;
        rom[70][21] = -8'd23;
        rom[70][22] = 8'd26;
        rom[70][23] = -8'd19;
        rom[70][24] = 8'd18;
        rom[70][25] = -8'd14;
        rom[70][26] = -8'd19;
        rom[70][27] = -8'd51;
        rom[70][28] = 8'd19;
        rom[70][29] = -8'd12;
        rom[70][30] = -8'd16;
        rom[70][31] = 8'd32;
        rom[71][0] = -8'd35;
        rom[71][1] = 8'd18;
        rom[71][2] = 8'd18;
        rom[71][3] = 8'd30;
        rom[71][4] = 8'd4;
        rom[71][5] = -8'd74;
        rom[71][6] = -8'd1;
        rom[71][7] = 8'd6;
        rom[71][8] = 8'd12;
        rom[71][9] = 8'd16;
        rom[71][10] = -8'd21;
        rom[71][11] = -8'd25;
        rom[71][12] = 8'd34;
        rom[71][13] = -8'd9;
        rom[71][14] = -8'd41;
        rom[71][15] = -8'd8;
        rom[71][16] = 8'd7;
        rom[71][17] = 8'd22;
        rom[71][18] = -8'd10;
        rom[71][19] = 8'd7;
        rom[71][20] = -8'd10;
        rom[71][21] = 8'd3;
        rom[71][22] = -8'd4;
        rom[71][23] = -8'd19;
        rom[71][24] = -8'd1;
        rom[71][25] = -8'd12;
        rom[71][26] = 8'd25;
        rom[71][27] = 8'd16;
        rom[71][28] = 8'd17;
        rom[71][29] = 8'd2;
        rom[71][30] = 8'd12;
        rom[71][31] = -8'd10;
        rom[72][0] = 8'd7;
        rom[72][1] = 8'd27;
        rom[72][2] = 8'd19;
        rom[72][3] = -8'd10;
        rom[72][4] = -8'd6;
        rom[72][5] = 8'd6;
        rom[72][6] = -8'd18;
        rom[72][7] = -8'd2;
        rom[72][8] = -8'd22;
        rom[72][9] = -8'd1;
        rom[72][10] = -8'd13;
        rom[72][11] = 8'd13;
        rom[72][12] = 8'd14;
        rom[72][13] = -8'd39;
        rom[72][14] = 8'd47;
        rom[72][15] = -8'd14;
        rom[72][16] = 8'd16;
        rom[72][17] = -8'd17;
        rom[72][18] = -8'd7;
        rom[72][19] = -8'd31;
        rom[72][20] = -8'd4;
        rom[72][21] = -8'd8;
        rom[72][22] = -8'd8;
        rom[72][23] = -8'd3;
        rom[72][24] = 8'd29;
        rom[72][25] = -8'd15;
        rom[72][26] = 8'd9;
        rom[72][27] = 8'd27;
        rom[72][28] = -8'd18;
        rom[72][29] = -8'd13;
        rom[72][30] = -8'd5;
        rom[72][31] = -8'd4;
        rom[73][0] = -8'd2;
        rom[73][1] = -8'd4;
        rom[73][2] = -8'd7;
        rom[73][3] = 8'd20;
        rom[73][4] = -8'd22;
        rom[73][5] = -8'd9;
        rom[73][6] = 8'd18;
        rom[73][7] = -8'd4;
        rom[73][8] = -8'd45;
        rom[73][9] = 8'd19;
        rom[73][10] = 8'd27;
        rom[73][11] = 8'd22;
        rom[73][12] = -8'd5;
        rom[73][13] = -8'd31;
        rom[73][14] = 8'd4;
        rom[73][15] = 8'd30;
        rom[73][16] = -8'd5;
        rom[73][17] = -8'd6;
        rom[73][18] = -8'd11;
        rom[73][19] = 8'd34;
        rom[73][20] = 8'd39;
        rom[73][21] = -8'd10;
        rom[73][22] = 8'd11;
        rom[73][23] = -8'd3;
        rom[73][24] = 8'd37;
        rom[73][25] = -8'd7;
        rom[73][26] = 8'd19;
        rom[73][27] = 8'd1;
        rom[73][28] = -8'd8;
        rom[73][29] = -8'd1;
        rom[73][30] = -8'd21;
        rom[73][31] = 8'd12;
        rom[74][0] = 8'd57;
        rom[74][1] = -8'd5;
        rom[74][2] = -8'd20;
        rom[74][3] = 8'd10;
        rom[74][4] = 8'd10;
        rom[74][5] = 8'd32;
        rom[74][6] = 8'd6;
        rom[74][7] = -8'd34;
        rom[74][8] = 8'd7;
        rom[74][9] = 8'd22;
        rom[74][10] = 8'd38;
        rom[74][11] = -8'd19;
        rom[74][12] = -8'd29;
        rom[74][13] = -8'd10;
        rom[74][14] = 8'd26;
        rom[74][15] = 8'd0;
        rom[74][16] = 8'd10;
        rom[74][17] = 8'd57;
        rom[74][18] = -8'd21;
        rom[74][19] = 8'd26;
        rom[74][20] = -8'd7;
        rom[74][21] = 8'd4;
        rom[74][22] = 8'd42;
        rom[74][23] = -8'd41;
        rom[74][24] = 8'd36;
        rom[74][25] = -8'd14;
        rom[74][26] = -8'd5;
        rom[74][27] = -8'd16;
        rom[74][28] = -8'd14;
        rom[74][29] = -8'd10;
        rom[74][30] = 8'd33;
        rom[74][31] = 8'd8;
        rom[75][0] = 8'd41;
        rom[75][1] = -8'd36;
        rom[75][2] = -8'd42;
        rom[75][3] = -8'd9;
        rom[75][4] = 8'd14;
        rom[75][5] = -8'd17;
        rom[75][6] = 8'd29;
        rom[75][7] = -8'd51;
        rom[75][8] = 8'd45;
        rom[75][9] = 8'd13;
        rom[75][10] = -8'd10;
        rom[75][11] = -8'd10;
        rom[75][12] = -8'd23;
        rom[75][13] = 8'd25;
        rom[75][14] = 8'd22;
        rom[75][15] = 8'd13;
        rom[75][16] = 8'd39;
        rom[75][17] = -8'd6;
        rom[75][18] = 8'd17;
        rom[75][19] = 8'd26;
        rom[75][20] = 8'd45;
        rom[75][21] = -8'd6;
        rom[75][22] = -8'd5;
        rom[75][23] = -8'd49;
        rom[75][24] = -8'd20;
        rom[75][25] = -8'd26;
        rom[75][26] = 8'd1;
        rom[75][27] = 8'd5;
        rom[75][28] = 8'd3;
        rom[75][29] = -8'd14;
        rom[75][30] = 8'd38;
        rom[75][31] = -8'd19;
        rom[76][0] = 8'd46;
        rom[76][1] = 8'd20;
        rom[76][2] = -8'd5;
        rom[76][3] = -8'd5;
        rom[76][4] = -8'd18;
        rom[76][5] = -8'd17;
        rom[76][6] = -8'd5;
        rom[76][7] = -8'd13;
        rom[76][8] = -8'd15;
        rom[76][9] = 8'd1;
        rom[76][10] = 8'd22;
        rom[76][11] = 8'd13;
        rom[76][12] = 8'd41;
        rom[76][13] = -8'd3;
        rom[76][14] = -8'd13;
        rom[76][15] = 8'd26;
        rom[76][16] = 8'd44;
        rom[76][17] = 8'd11;
        rom[76][18] = 8'd0;
        rom[76][19] = -8'd3;
        rom[76][20] = 8'd37;
        rom[76][21] = 8'd13;
        rom[76][22] = -8'd25;
        rom[76][23] = 8'd32;
        rom[76][24] = -8'd1;
        rom[76][25] = 8'd30;
        rom[76][26] = 8'd16;
        rom[76][27] = 8'd52;
        rom[76][28] = -8'd28;
        rom[76][29] = -8'd1;
        rom[76][30] = -8'd75;
        rom[76][31] = 8'd16;
        rom[77][0] = -8'd41;
        rom[77][1] = -8'd29;
        rom[77][2] = -8'd11;
        rom[77][3] = 8'd4;
        rom[77][4] = 8'd21;
        rom[77][5] = -8'd16;
        rom[77][6] = -8'd5;
        rom[77][7] = -8'd30;
        rom[77][8] = -8'd30;
        rom[77][9] = -8'd48;
        rom[77][10] = 8'd7;
        rom[77][11] = -8'd3;
        rom[77][12] = -8'd7;
        rom[77][13] = -8'd35;
        rom[77][14] = -8'd4;
        rom[77][15] = 8'd48;
        rom[77][16] = -8'd23;
        rom[77][17] = -8'd21;
        rom[77][18] = 8'd21;
        rom[77][19] = 8'd6;
        rom[77][20] = 8'd5;
        rom[77][21] = -8'd24;
        rom[77][22] = -8'd33;
        rom[77][23] = 8'd24;
        rom[77][24] = -8'd1;
        rom[77][25] = -8'd11;
        rom[77][26] = -8'd8;
        rom[77][27] = 8'd43;
        rom[77][28] = -8'd20;
        rom[77][29] = -8'd5;
        rom[77][30] = -8'd26;
        rom[77][31] = -8'd47;
        rom[78][0] = -8'd60;
        rom[78][1] = 8'd19;
        rom[78][2] = 8'd55;
        rom[78][3] = 8'd19;
        rom[78][4] = 8'd20;
        rom[78][5] = -8'd95;
        rom[78][6] = 8'd2;
        rom[78][7] = 8'd14;
        rom[78][8] = 8'd21;
        rom[78][9] = 8'd10;
        rom[78][10] = 8'd6;
        rom[78][11] = -8'd7;
        rom[78][12] = 8'd3;
        rom[78][13] = -8'd23;
        rom[78][14] = -8'd3;
        rom[78][15] = 8'd14;
        rom[78][16] = -8'd15;
        rom[78][17] = -8'd29;
        rom[78][18] = 8'd10;
        rom[78][19] = 8'd15;
        rom[78][20] = 8'd9;
        rom[78][21] = -8'd17;
        rom[78][22] = -8'd29;
        rom[78][23] = 8'd29;
        rom[78][24] = 8'd7;
        rom[78][25] = 8'd62;
        rom[78][26] = -8'd19;
        rom[78][27] = 8'd7;
        rom[78][28] = -8'd2;
        rom[78][29] = -8'd8;
        rom[78][30] = -8'd9;
        rom[78][31] = -8'd13;
        rom[79][0] = -8'd14;
        rom[79][1] = 8'd30;
        rom[79][2] = 8'd28;
        rom[79][3] = 8'd3;
        rom[79][4] = 8'd12;
        rom[79][5] = -8'd34;
        rom[79][6] = 8'd31;
        rom[79][7] = -8'd9;
        rom[79][8] = -8'd18;
        rom[79][9] = 8'd24;
        rom[79][10] = -8'd47;
        rom[79][11] = -8'd21;
        rom[79][12] = -8'd38;
        rom[79][13] = -8'd8;
        rom[79][14] = -8'd12;
        rom[79][15] = 8'd13;
        rom[79][16] = -8'd16;
        rom[79][17] = 8'd8;
        rom[79][18] = 8'd24;
        rom[79][19] = 8'd13;
        rom[79][20] = 8'd15;
        rom[79][21] = -8'd7;
        rom[79][22] = 8'd3;
        rom[79][23] = -8'd17;
        rom[79][24] = 8'd9;
        rom[79][25] = -8'd16;
        rom[79][26] = -8'd9;
        rom[79][27] = 8'd12;
        rom[79][28] = -8'd2;
        rom[79][29] = -8'd12;
        rom[79][30] = -8'd11;
        rom[79][31] = 8'd14;
        rom[80][0] = 8'd26;
        rom[80][1] = 8'd31;
        rom[80][2] = -8'd27;
        rom[80][3] = 8'd5;
        rom[80][4] = -8'd4;
        rom[80][5] = 8'd26;
        rom[80][6] = -8'd39;
        rom[80][7] = -8'd11;
        rom[80][8] = -8'd3;
        rom[80][9] = 8'd11;
        rom[80][10] = -8'd8;
        rom[80][11] = -8'd7;
        rom[80][12] = 8'd39;
        rom[80][13] = 8'd7;
        rom[80][14] = -8'd17;
        rom[80][15] = -8'd19;
        rom[80][16] = 8'd47;
        rom[80][17] = -8'd35;
        rom[80][18] = 8'd12;
        rom[80][19] = -8'd41;
        rom[80][20] = 8'd6;
        rom[80][21] = -8'd27;
        rom[80][22] = 8'd0;
        rom[80][23] = 8'd1;
        rom[80][24] = 8'd7;
        rom[80][25] = 8'd11;
        rom[80][26] = 8'd5;
        rom[80][27] = 8'd10;
        rom[80][28] = -8'd28;
        rom[80][29] = -8'd15;
        rom[80][30] = 8'd32;
        rom[80][31] = -8'd18;
        rom[81][0] = -8'd13;
        rom[81][1] = -8'd48;
        rom[81][2] = -8'd38;
        rom[81][3] = 8'd31;
        rom[81][4] = -8'd7;
        rom[81][5] = -8'd62;
        rom[81][6] = -8'd11;
        rom[81][7] = 8'd20;
        rom[81][8] = -8'd28;
        rom[81][9] = 8'd22;
        rom[81][10] = -8'd6;
        rom[81][11] = 8'd3;
        rom[81][12] = -8'd19;
        rom[81][13] = 8'd20;
        rom[81][14] = -8'd25;
        rom[81][15] = -8'd20;
        rom[81][16] = -8'd53;
        rom[81][17] = 8'd18;
        rom[81][18] = -8'd5;
        rom[81][19] = 8'd16;
        rom[81][20] = 8'd17;
        rom[81][21] = -8'd4;
        rom[81][22] = 8'd3;
        rom[81][23] = 8'd24;
        rom[81][24] = 8'd19;
        rom[81][25] = -8'd3;
        rom[81][26] = -8'd13;
        rom[81][27] = 8'd25;
        rom[81][28] = -8'd1;
        rom[81][29] = 8'd3;
        rom[81][30] = -8'd23;
        rom[81][31] = 8'd4;
        rom[82][0] = 8'd10;
        rom[82][1] = -8'd33;
        rom[82][2] = -8'd8;
        rom[82][3] = 8'd23;
        rom[82][4] = 8'd28;
        rom[82][5] = -8'd14;
        rom[82][6] = -8'd10;
        rom[82][7] = 8'd50;
        rom[82][8] = -8'd25;
        rom[82][9] = -8'd37;
        rom[82][10] = 8'd5;
        rom[82][11] = -8'd11;
        rom[82][12] = -8'd30;
        rom[82][13] = -8'd16;
        rom[82][14] = -8'd14;
        rom[82][15] = -8'd34;
        rom[82][16] = -8'd78;
        rom[82][17] = -8'd33;
        rom[82][18] = -8'd23;
        rom[82][19] = -8'd17;
        rom[82][20] = 8'd27;
        rom[82][21] = -8'd14;
        rom[82][22] = 8'd9;
        rom[82][23] = 8'd24;
        rom[82][24] = -8'd2;
        rom[82][25] = 8'd40;
        rom[82][26] = -8'd52;
        rom[82][27] = -8'd14;
        rom[82][28] = 8'd6;
        rom[82][29] = 8'd3;
        rom[82][30] = 8'd3;
        rom[82][31] = 8'd1;
        rom[83][0] = -8'd15;
        rom[83][1] = -8'd18;
        rom[83][2] = 8'd11;
        rom[83][3] = -8'd20;
        rom[83][4] = -8'd15;
        rom[83][5] = 8'd24;
        rom[83][6] = -8'd11;
        rom[83][7] = -8'd26;
        rom[83][8] = -8'd12;
        rom[83][9] = -8'd27;
        rom[83][10] = 8'd35;
        rom[83][11] = 8'd12;
        rom[83][12] = -8'd7;
        rom[83][13] = -8'd16;
        rom[83][14] = -8'd4;
        rom[83][15] = 8'd22;
        rom[83][16] = 8'd10;
        rom[83][17] = 8'd0;
        rom[83][18] = 8'd11;
        rom[83][19] = 8'd17;
        rom[83][20] = 8'd45;
        rom[83][21] = -8'd5;
        rom[83][22] = -8'd12;
        rom[83][23] = 8'd13;
        rom[83][24] = 8'd2;
        rom[83][25] = 8'd22;
        rom[83][26] = -8'd4;
        rom[83][27] = 8'd0;
        rom[83][28] = 8'd12;
        rom[83][29] = -8'd12;
        rom[83][30] = -8'd23;
        rom[83][31] = -8'd26;
        rom[84][0] = -8'd10;
        rom[84][1] = 8'd27;
        rom[84][2] = -8'd21;
        rom[84][3] = 8'd45;
        rom[84][4] = -8'd13;
        rom[84][5] = 8'd13;
        rom[84][6] = 8'd22;
        rom[84][7] = -8'd36;
        rom[84][8] = 8'd8;
        rom[84][9] = 8'd17;
        rom[84][10] = 8'd12;
        rom[84][11] = -8'd31;
        rom[84][12] = -8'd1;
        rom[84][13] = 8'd5;
        rom[84][14] = -8'd28;
        rom[84][15] = 8'd5;
        rom[84][16] = -8'd3;
        rom[84][17] = 8'd12;
        rom[84][18] = -8'd9;
        rom[84][19] = -8'd9;
        rom[84][20] = 8'd4;
        rom[84][21] = -8'd7;
        rom[84][22] = -8'd31;
        rom[84][23] = -8'd12;
        rom[84][24] = -8'd27;
        rom[84][25] = 8'd2;
        rom[84][26] = 8'd1;
        rom[84][27] = 8'd12;
        rom[84][28] = -8'd9;
        rom[84][29] = -8'd6;
        rom[84][30] = -8'd35;
        rom[84][31] = -8'd26;
        rom[85][0] = 8'd12;
        rom[85][1] = -8'd53;
        rom[85][2] = 8'd24;
        rom[85][3] = 8'd5;
        rom[85][4] = -8'd13;
        rom[85][5] = -8'd89;
        rom[85][6] = 8'd10;
        rom[85][7] = -8'd4;
        rom[85][8] = 8'd19;
        rom[85][9] = -8'd29;
        rom[85][10] = -8'd11;
        rom[85][11] = 8'd31;
        rom[85][12] = 8'd17;
        rom[85][13] = -8'd14;
        rom[85][14] = 8'd6;
        rom[85][15] = 8'd24;
        rom[85][16] = -8'd12;
        rom[85][17] = -8'd9;
        rom[85][18] = 8'd3;
        rom[85][19] = 8'd9;
        rom[85][20] = -8'd28;
        rom[85][21] = -8'd19;
        rom[85][22] = 8'd14;
        rom[85][23] = -8'd1;
        rom[85][24] = -8'd28;
        rom[85][25] = -8'd64;
        rom[85][26] = -8'd33;
        rom[85][27] = 8'd9;
        rom[85][28] = -8'd42;
        rom[85][29] = 8'd9;
        rom[85][30] = 8'd53;
        rom[85][31] = -8'd8;
        rom[86][0] = -8'd99;
        rom[86][1] = -8'd25;
        rom[86][2] = -8'd6;
        rom[86][3] = 8'd2;
        rom[86][4] = -8'd35;
        rom[86][5] = -8'd37;
        rom[86][6] = -8'd7;
        rom[86][7] = 8'd37;
        rom[86][8] = 8'd10;
        rom[86][9] = 8'd29;
        rom[86][10] = 8'd17;
        rom[86][11] = 8'd2;
        rom[86][12] = -8'd5;
        rom[86][13] = -8'd21;
        rom[86][14] = -8'd27;
        rom[86][15] = -8'd16;
        rom[86][16] = -8'd6;
        rom[86][17] = 8'd37;
        rom[86][18] = -8'd18;
        rom[86][19] = -8'd11;
        rom[86][20] = 8'd39;
        rom[86][21] = 8'd13;
        rom[86][22] = 8'd15;
        rom[86][23] = 8'd8;
        rom[86][24] = 8'd16;
        rom[86][25] = 8'd12;
        rom[86][26] = -8'd28;
        rom[86][27] = 8'd17;
        rom[86][28] = 8'd15;
        rom[86][29] = -8'd12;
        rom[86][30] = 8'd14;
        rom[86][31] = -8'd2;
        rom[87][0] = 8'd12;
        rom[87][1] = 8'd26;
        rom[87][2] = 8'd19;
        rom[87][3] = 8'd21;
        rom[87][4] = -8'd4;
        rom[87][5] = -8'd53;
        rom[87][6] = -8'd19;
        rom[87][7] = 8'd18;
        rom[87][8] = 8'd35;
        rom[87][9] = -8'd4;
        rom[87][10] = 8'd22;
        rom[87][11] = -8'd2;
        rom[87][12] = 8'd20;
        rom[87][13] = 8'd11;
        rom[87][14] = -8'd33;
        rom[87][15] = 8'd8;
        rom[87][16] = -8'd32;
        rom[87][17] = 8'd21;
        rom[87][18] = 8'd13;
        rom[87][19] = 8'd25;
        rom[87][20] = -8'd18;
        rom[87][21] = 8'd11;
        rom[87][22] = 8'd8;
        rom[87][23] = -8'd23;
        rom[87][24] = 8'd8;
        rom[87][25] = -8'd32;
        rom[87][26] = 8'd10;
        rom[87][27] = 8'd23;
        rom[87][28] = 8'd23;
        rom[87][29] = 8'd4;
        rom[87][30] = 8'd0;
        rom[87][31] = 8'd5;
        rom[88][0] = 8'd7;
        rom[88][1] = -8'd38;
        rom[88][2] = -8'd24;
        rom[88][3] = -8'd63;
        rom[88][4] = 8'd30;
        rom[88][5] = 8'd5;
        rom[88][6] = 8'd16;
        rom[88][7] = -8'd14;
        rom[88][8] = -8'd22;
        rom[88][9] = -8'd11;
        rom[88][10] = 8'd21;
        rom[88][11] = 8'd31;
        rom[88][12] = 8'd24;
        rom[88][13] = 8'd33;
        rom[88][14] = 8'd18;
        rom[88][15] = 8'd7;
        rom[88][16] = 8'd1;
        rom[88][17] = -8'd62;
        rom[88][18] = -8'd9;
        rom[88][19] = 8'd7;
        rom[88][20] = -8'd8;
        rom[88][21] = -8'd70;
        rom[88][22] = -8'd15;
        rom[88][23] = 8'd0;
        rom[88][24] = 8'd5;
        rom[88][25] = -8'd1;
        rom[88][26] = -8'd26;
        rom[88][27] = -8'd15;
        rom[88][28] = -8'd45;
        rom[88][29] = -8'd8;
        rom[88][30] = 8'd34;
        rom[88][31] = -8'd25;
        rom[89][0] = -8'd6;
        rom[89][1] = -8'd35;
        rom[89][2] = 8'd10;
        rom[89][3] = -8'd10;
        rom[89][4] = -8'd19;
        rom[89][5] = -8'd41;
        rom[89][6] = 8'd8;
        rom[89][7] = 8'd8;
        rom[89][8] = 8'd12;
        rom[89][9] = 8'd12;
        rom[89][10] = -8'd32;
        rom[89][11] = -8'd16;
        rom[89][12] = -8'd48;
        rom[89][13] = 8'd24;
        rom[89][14] = 8'd9;
        rom[89][15] = -8'd32;
        rom[89][16] = -8'd14;
        rom[89][17] = -8'd4;
        rom[89][18] = 8'd31;
        rom[89][19] = 8'd11;
        rom[89][20] = -8'd35;
        rom[89][21] = 8'd1;
        rom[89][22] = 8'd3;
        rom[89][23] = -8'd53;
        rom[89][24] = 8'd15;
        rom[89][25] = -8'd33;
        rom[89][26] = -8'd11;
        rom[89][27] = -8'd4;
        rom[89][28] = -8'd11;
        rom[89][29] = -8'd17;
        rom[89][30] = 8'd2;
        rom[89][31] = -8'd27;
        rom[90][0] = 8'd14;
        rom[90][1] = 8'd2;
        rom[90][2] = -8'd64;
        rom[90][3] = 8'd3;
        rom[90][4] = 8'd19;
        rom[90][5] = 8'd10;
        rom[90][6] = 8'd2;
        rom[90][7] = 8'd8;
        rom[90][8] = -8'd11;
        rom[90][9] = 8'd27;
        rom[90][10] = -8'd15;
        rom[90][11] = 8'd24;
        rom[90][12] = 8'd10;
        rom[90][13] = -8'd8;
        rom[90][14] = -8'd21;
        rom[90][15] = -8'd7;
        rom[90][16] = -8'd24;
        rom[90][17] = -8'd20;
        rom[90][18] = -8'd2;
        rom[90][19] = 8'd6;
        rom[90][20] = -8'd1;
        rom[90][21] = 8'd9;
        rom[90][22] = 8'd13;
        rom[90][23] = 8'd7;
        rom[90][24] = 8'd23;
        rom[90][25] = -8'd23;
        rom[90][26] = 8'd10;
        rom[90][27] = -8'd2;
        rom[90][28] = 8'd17;
        rom[90][29] = 8'd2;
        rom[90][30] = -8'd24;
        rom[90][31] = 8'd16;
        rom[91][0] = -8'd14;
        rom[91][1] = 8'd6;
        rom[91][2] = 8'd26;
        rom[91][3] = -8'd3;
        rom[91][4] = 8'd17;
        rom[91][5] = -8'd26;
        rom[91][6] = 8'd35;
        rom[91][7] = -8'd31;
        rom[91][8] = -8'd12;
        rom[91][9] = 8'd0;
        rom[91][10] = 8'd8;
        rom[91][11] = 8'd3;
        rom[91][12] = 8'd17;
        rom[91][13] = -8'd12;
        rom[91][14] = 8'd7;
        rom[91][15] = 8'd7;
        rom[91][16] = -8'd3;
        rom[91][17] = -8'd6;
        rom[91][18] = 8'd17;
        rom[91][19] = 8'd2;
        rom[91][20] = 8'd3;
        rom[91][21] = -8'd9;
        rom[91][22] = -8'd2;
        rom[91][23] = 8'd22;
        rom[91][24] = -8'd7;
        rom[91][25] = -8'd10;
        rom[91][26] = 8'd10;
        rom[91][27] = -8'd11;
        rom[91][28] = 8'd25;
        rom[91][29] = -8'd17;
        rom[91][30] = 8'd7;
        rom[91][31] = 8'd5;
        rom[92][0] = -8'd5;
        rom[92][1] = 8'd15;
        rom[92][2] = 8'd1;
        rom[92][3] = 8'd64;
        rom[92][4] = 8'd17;
        rom[92][5] = 8'd17;
        rom[92][6] = 8'd6;
        rom[92][7] = -8'd1;
        rom[92][8] = -8'd22;
        rom[92][9] = 8'd10;
        rom[92][10] = 8'd5;
        rom[92][11] = 8'd5;
        rom[92][12] = -8'd28;
        rom[92][13] = -8'd27;
        rom[92][14] = 8'd12;
        rom[92][15] = -8'd14;
        rom[92][16] = -8'd7;
        rom[92][17] = -8'd9;
        rom[92][18] = 8'd9;
        rom[92][19] = 8'd0;
        rom[92][20] = -8'd12;
        rom[92][21] = -8'd7;
        rom[92][22] = -8'd1;
        rom[92][23] = -8'd1;
        rom[92][24] = -8'd22;
        rom[92][25] = 8'd10;
        rom[92][26] = 8'd21;
        rom[92][27] = 8'd33;
        rom[92][28] = -8'd7;
        rom[92][29] = -8'd11;
        rom[92][30] = -8'd8;
        rom[92][31] = -8'd16;
        rom[93][0] = -8'd44;
        rom[93][1] = -8'd27;
        rom[93][2] = 8'd33;
        rom[93][3] = -8'd29;
        rom[93][4] = 8'd14;
        rom[93][5] = -8'd20;
        rom[93][6] = 8'd18;
        rom[93][7] = -8'd9;
        rom[93][8] = 8'd31;
        rom[93][9] = 8'd45;
        rom[93][10] = 8'd23;
        rom[93][11] = -8'd23;
        rom[93][12] = 8'd4;
        rom[93][13] = 8'd34;
        rom[93][14] = 8'd17;
        rom[93][15] = 8'd21;
        rom[93][16] = 8'd18;
        rom[93][17] = 8'd26;
        rom[93][18] = -8'd37;
        rom[93][19] = 8'd39;
        rom[93][20] = -8'd11;
        rom[93][21] = 8'd13;
        rom[93][22] = -8'd42;
        rom[93][23] = -8'd21;
        rom[93][24] = -8'd40;
        rom[93][25] = 8'd2;
        rom[93][26] = 8'd10;
        rom[93][27] = 8'd12;
        rom[93][28] = 8'd44;
        rom[93][29] = 8'd9;
        rom[93][30] = 8'd16;
        rom[93][31] = -8'd51;
        rom[94][0] = -8'd20;
        rom[94][1] = 8'd54;
        rom[94][2] = -8'd27;
        rom[94][3] = -8'd14;
        rom[94][4] = -8'd13;
        rom[94][5] = -8'd20;
        rom[94][6] = -8'd10;
        rom[94][7] = -8'd50;
        rom[94][8] = 8'd7;
        rom[94][9] = -8'd3;
        rom[94][10] = -8'd24;
        rom[94][11] = -8'd56;
        rom[94][12] = -8'd16;
        rom[94][13] = 8'd15;
        rom[94][14] = 8'd13;
        rom[94][15] = -8'd15;
        rom[94][16] = 8'd27;
        rom[94][17] = 8'd27;
        rom[94][18] = -8'd9;
        rom[94][19] = -8'd13;
        rom[94][20] = -8'd17;
        rom[94][21] = 8'd16;
        rom[94][22] = -8'd38;
        rom[94][23] = -8'd16;
        rom[94][24] = 8'd14;
        rom[94][25] = 8'd4;
        rom[94][26] = -8'd15;
        rom[94][27] = -8'd7;
        rom[94][28] = 8'd8;
        rom[94][29] = 8'd4;
        rom[94][30] = 8'd2;
        rom[94][31] = -8'd14;
        rom[95][0] = 8'd32;
        rom[95][1] = -8'd2;
        rom[95][2] = -8'd51;
        rom[95][3] = 8'd6;
        rom[95][4] = 8'd28;
        rom[95][5] = 8'd65;
        rom[95][6] = 8'd2;
        rom[95][7] = -8'd38;
        rom[95][8] = -8'd43;
        rom[95][9] = -8'd53;
        rom[95][10] = -8'd33;
        rom[95][11] = -8'd16;
        rom[95][12] = -8'd18;
        rom[95][13] = -8'd12;
        rom[95][14] = -8'd29;
        rom[95][15] = 8'd4;
        rom[95][16] = -8'd29;
        rom[95][17] = -8'd33;
        rom[95][18] = -8'd14;
        rom[95][19] = -8'd21;
        rom[95][20] = -8'd7;
        rom[95][21] = -8'd38;
        rom[95][22] = 8'd67;
        rom[95][23] = -8'd7;
        rom[95][24] = 8'd17;
        rom[95][25] = 8'd23;
        rom[95][26] = -8'd16;
        rom[95][27] = -8'd46;
        rom[95][28] = -8'd2;
        rom[95][29] = -8'd4;
        rom[95][30] = 8'd3;
        rom[95][31] = 8'd13;
        rom[96][0] = -8'd40;
        rom[96][1] = 8'd22;
        rom[96][2] = -8'd1;
        rom[96][3] = -8'd8;
        rom[96][4] = 8'd30;
        rom[96][5] = -8'd25;
        rom[96][6] = 8'd20;
        rom[96][7] = 8'd2;
        rom[96][8] = 8'd15;
        rom[96][9] = -8'd12;
        rom[96][10] = -8'd22;
        rom[96][11] = -8'd29;
        rom[96][12] = -8'd25;
        rom[96][13] = -8'd9;
        rom[96][14] = 8'd1;
        rom[96][15] = -8'd9;
        rom[96][16] = 8'd12;
        rom[96][17] = 8'd14;
        rom[96][18] = -8'd4;
        rom[96][19] = 8'd16;
        rom[96][20] = -8'd7;
        rom[96][21] = 8'd48;
        rom[96][22] = -8'd5;
        rom[96][23] = 8'd10;
        rom[96][24] = -8'd14;
        rom[96][25] = 8'd22;
        rom[96][26] = 8'd1;
        rom[96][27] = -8'd10;
        rom[96][28] = 8'd4;
        rom[96][29] = -8'd2;
        rom[96][30] = -8'd3;
        rom[96][31] = 8'd1;
        rom[97][0] = 8'd17;
        rom[97][1] = -8'd18;
        rom[97][2] = -8'd36;
        rom[97][3] = -8'd13;
        rom[97][4] = -8'd24;
        rom[97][5] = 8'd20;
        rom[97][6] = -8'd32;
        rom[97][7] = -8'd48;
        rom[97][8] = -8'd19;
        rom[97][9] = -8'd5;
        rom[97][10] = -8'd24;
        rom[97][11] = -8'd19;
        rom[97][12] = -8'd18;
        rom[97][13] = 8'd15;
        rom[97][14] = -8'd30;
        rom[97][15] = -8'd10;
        rom[97][16] = 8'd10;
        rom[97][17] = -8'd37;
        rom[97][18] = 8'd0;
        rom[97][19] = -8'd3;
        rom[97][20] = 8'd20;
        rom[97][21] = -8'd2;
        rom[97][22] = -8'd33;
        rom[97][23] = 8'd31;
        rom[97][24] = 8'd31;
        rom[97][25] = -8'd19;
        rom[97][26] = -8'd3;
        rom[97][27] = -8'd20;
        rom[97][28] = 8'd8;
        rom[97][29] = -8'd2;
        rom[97][30] = -8'd14;
        rom[97][31] = -8'd2;
        rom[98][0] = -8'd65;
        rom[98][1] = -8'd3;
        rom[98][2] = 8'd29;
        rom[98][3] = -8'd11;
        rom[98][4] = -8'd4;
        rom[98][5] = 8'd39;
        rom[98][6] = 8'd6;
        rom[98][7] = -8'd12;
        rom[98][8] = 8'd45;
        rom[98][9] = -8'd55;
        rom[98][10] = -8'd43;
        rom[98][11] = -8'd56;
        rom[98][12] = -8'd11;
        rom[98][13] = -8'd18;
        rom[98][14] = 8'd12;
        rom[98][15] = -8'd26;
        rom[98][16] = 8'd35;
        rom[98][17] = 8'd16;
        rom[98][18] = 8'd22;
        rom[98][19] = -8'd48;
        rom[98][20] = -8'd18;
        rom[98][21] = -8'd29;
        rom[98][22] = 8'd40;
        rom[98][23] = -8'd55;
        rom[98][24] = -8'd25;
        rom[98][25] = -8'd33;
        rom[98][26] = -8'd10;
        rom[98][27] = -8'd27;
        rom[98][28] = 8'd12;
        rom[98][29] = -8'd16;
        rom[98][30] = -8'd26;
        rom[98][31] = 8'd4;
        rom[99][0] = -8'd31;
        rom[99][1] = -8'd9;
        rom[99][2] = 8'd3;
        rom[99][3] = 8'd25;
        rom[99][4] = -8'd28;
        rom[99][5] = -8'd12;
        rom[99][6] = 8'd28;
        rom[99][7] = -8'd27;
        rom[99][8] = 8'd13;
        rom[99][9] = -8'd25;
        rom[99][10] = 8'd14;
        rom[99][11] = 8'd22;
        rom[99][12] = -8'd34;
        rom[99][13] = 8'd12;
        rom[99][14] = -8'd5;
        rom[99][15] = -8'd76;
        rom[99][16] = 8'd16;
        rom[99][17] = -8'd37;
        rom[99][18] = 8'd2;
        rom[99][19] = -8'd15;
        rom[99][20] = -8'd32;
        rom[99][21] = 8'd7;
        rom[99][22] = 8'd22;
        rom[99][23] = -8'd29;
        rom[99][24] = 8'd28;
        rom[99][25] = -8'd25;
        rom[99][26] = 8'd16;
        rom[99][27] = -8'd23;
        rom[99][28] = -8'd1;
        rom[99][29] = 8'd4;
        rom[99][30] = 8'd34;
        rom[99][31] = 8'd9;
        rom[100][0] = -8'd3;
        rom[100][1] = -8'd30;
        rom[100][2] = -8'd37;
        rom[100][3] = -8'd1;
        rom[100][4] = 8'd7;
        rom[100][5] = 8'd11;
        rom[100][6] = -8'd14;
        rom[100][7] = -8'd13;
        rom[100][8] = -8'd8;
        rom[100][9] = -8'd3;
        rom[100][10] = 8'd35;
        rom[100][11] = 8'd44;
        rom[100][12] = 8'd24;
        rom[100][13] = 8'd22;
        rom[100][14] = -8'd54;
        rom[100][15] = 8'd44;
        rom[100][16] = 8'd1;
        rom[100][17] = 8'd32;
        rom[100][18] = 8'd6;
        rom[100][19] = -8'd49;
        rom[100][20] = 8'd20;
        rom[100][21] = -8'd26;
        rom[100][22] = -8'd36;
        rom[100][23] = 8'd47;
        rom[100][24] = 8'd28;
        rom[100][25] = 8'd3;
        rom[100][26] = -8'd43;
        rom[100][27] = -8'd38;
        rom[100][28] = 8'd11;
        rom[100][29] = 8'd0;
        rom[100][30] = 8'd8;
        rom[100][31] = 8'd33;
        rom[101][0] = -8'd78;
        rom[101][1] = 8'd21;
        rom[101][2] = 8'd11;
        rom[101][3] = -8'd15;
        rom[101][4] = -8'd97;
        rom[101][5] = 8'd38;
        rom[101][6] = 8'd10;
        rom[101][7] = 8'd7;
        rom[101][8] = 8'd46;
        rom[101][9] = -8'd34;
        rom[101][10] = 8'd25;
        rom[101][11] = -8'd15;
        rom[101][12] = -8'd96;
        rom[101][13] = 8'd41;
        rom[101][14] = 8'd23;
        rom[101][15] = -8'd28;
        rom[101][16] = -8'd9;
        rom[101][17] = -8'd1;
        rom[101][18] = -8'd8;
        rom[101][19] = 8'd17;
        rom[101][20] = 8'd28;
        rom[101][21] = -8'd2;
        rom[101][22] = 8'd3;
        rom[101][23] = -8'd27;
        rom[101][24] = -8'd69;
        rom[101][25] = 8'd39;
        rom[101][26] = -8'd23;
        rom[101][27] = -8'd31;
        rom[101][28] = -8'd1;
        rom[101][29] = 8'd5;
        rom[101][30] = -8'd12;
        rom[101][31] = -8'd6;
        rom[102][0] = -8'd14;
        rom[102][1] = 8'd14;
        rom[102][2] = -8'd6;
        rom[102][3] = -8'd43;
        rom[102][4] = 8'd9;
        rom[102][5] = 8'd35;
        rom[102][6] = -8'd9;
        rom[102][7] = 8'd5;
        rom[102][8] = 8'd23;
        rom[102][9] = -8'd32;
        rom[102][10] = -8'd11;
        rom[102][11] = 8'd19;
        rom[102][12] = -8'd28;
        rom[102][13] = -8'd7;
        rom[102][14] = 8'd6;
        rom[102][15] = 8'd4;
        rom[102][16] = -8'd4;
        rom[102][17] = 8'd45;
        rom[102][18] = -8'd41;
        rom[102][19] = -8'd10;
        rom[102][20] = -8'd5;
        rom[102][21] = -8'd17;
        rom[102][22] = 8'd26;
        rom[102][23] = 8'd12;
        rom[102][24] = 8'd16;
        rom[102][25] = -8'd36;
        rom[102][26] = -8'd5;
        rom[102][27] = -8'd6;
        rom[102][28] = 8'd16;
        rom[102][29] = -8'd10;
        rom[102][30] = -8'd33;
        rom[102][31] = 8'd25;
        rom[103][0] = -8'd12;
        rom[103][1] = 8'd9;
        rom[103][2] = 8'd0;
        rom[103][3] = -8'd7;
        rom[103][4] = 8'd16;
        rom[103][5] = -8'd33;
        rom[103][6] = -8'd23;
        rom[103][7] = 8'd12;
        rom[103][8] = -8'd33;
        rom[103][9] = 8'd12;
        rom[103][10] = 8'd26;
        rom[103][11] = 8'd23;
        rom[103][12] = 8'd17;
        rom[103][13] = 8'd13;
        rom[103][14] = -8'd31;
        rom[103][15] = -8'd11;
        rom[103][16] = 8'd0;
        rom[103][17] = 8'd4;
        rom[103][18] = 8'd4;
        rom[103][19] = -8'd20;
        rom[103][20] = -8'd9;
        rom[103][21] = -8'd6;
        rom[103][22] = -8'd24;
        rom[103][23] = 8'd7;
        rom[103][24] = -8'd12;
        rom[103][25] = 8'd0;
        rom[103][26] = 8'd38;
        rom[103][27] = 8'd16;
        rom[103][28] = 8'd11;
        rom[103][29] = 8'd1;
        rom[103][30] = -8'd7;
        rom[103][31] = 8'd10;
        rom[104][0] = -8'd15;
        rom[104][1] = 8'd11;
        rom[104][2] = -8'd7;
        rom[104][3] = 8'd24;
        rom[104][4] = 8'd13;
        rom[104][5] = 8'd11;
        rom[104][6] = 8'd30;
        rom[104][7] = 8'd12;
        rom[104][8] = -8'd23;
        rom[104][9] = 8'd19;
        rom[104][10] = 8'd22;
        rom[104][11] = 8'd30;
        rom[104][12] = 8'd0;
        rom[104][13] = -8'd9;
        rom[104][14] = -8'd52;
        rom[104][15] = 8'd7;
        rom[104][16] = 8'd7;
        rom[104][17] = -8'd43;
        rom[104][18] = 8'd18;
        rom[104][19] = -8'd42;
        rom[104][20] = 8'd34;
        rom[104][21] = 8'd4;
        rom[104][22] = 8'd24;
        rom[104][23] = 8'd0;
        rom[104][24] = 8'd16;
        rom[104][25] = -8'd7;
        rom[104][26] = 8'd1;
        rom[104][27] = 8'd4;
        rom[104][28] = -8'd10;
        rom[104][29] = -8'd5;
        rom[104][30] = -8'd5;
        rom[104][31] = -8'd20;
        rom[105][0] = -8'd15;
        rom[105][1] = -8'd2;
        rom[105][2] = -8'd3;
        rom[105][3] = 8'd5;
        rom[105][4] = 8'd18;
        rom[105][5] = 8'd32;
        rom[105][6] = -8'd3;
        rom[105][7] = 8'd23;
        rom[105][8] = 8'd48;
        rom[105][9] = -8'd9;
        rom[105][10] = -8'd10;
        rom[105][11] = 8'd32;
        rom[105][12] = -8'd6;
        rom[105][13] = -8'd11;
        rom[105][14] = 8'd36;
        rom[105][15] = -8'd16;
        rom[105][16] = -8'd34;
        rom[105][17] = 8'd31;
        rom[105][18] = 8'd2;
        rom[105][19] = -8'd31;
        rom[105][20] = -8'd15;
        rom[105][21] = 8'd22;
        rom[105][22] = 8'd46;
        rom[105][23] = -8'd31;
        rom[105][24] = 8'd6;
        rom[105][25] = -8'd3;
        rom[105][26] = -8'd18;
        rom[105][27] = -8'd41;
        rom[105][28] = 8'd2;
        rom[105][29] = -8'd1;
        rom[105][30] = 8'd50;
        rom[105][31] = -8'd32;
        rom[106][0] = -8'd52;
        rom[106][1] = -8'd27;
        rom[106][2] = -8'd1;
        rom[106][3] = -8'd23;
        rom[106][4] = -8'd28;
        rom[106][5] = 8'd5;
        rom[106][6] = 8'd10;
        rom[106][7] = 8'd40;
        rom[106][8] = -8'd29;
        rom[106][9] = 8'd3;
        rom[106][10] = 8'd7;
        rom[106][11] = 8'd53;
        rom[106][12] = -8'd1;
        rom[106][13] = -8'd30;
        rom[106][14] = 8'd33;
        rom[106][15] = 8'd2;
        rom[106][16] = 8'd28;
        rom[106][17] = 8'd17;
        rom[106][18] = 8'd19;
        rom[106][19] = -8'd22;
        rom[106][20] = 8'd11;
        rom[106][21] = 8'd45;
        rom[106][22] = -8'd14;
        rom[106][23] = -8'd13;
        rom[106][24] = 8'd11;
        rom[106][25] = 8'd22;
        rom[106][26] = 8'd15;
        rom[106][27] = -8'd23;
        rom[106][28] = 8'd17;
        rom[106][29] = 8'd2;
        rom[106][30] = 8'd2;
        rom[106][31] = -8'd27;
        rom[107][0] = 8'd35;
        rom[107][1] = -8'd23;
        rom[107][2] = -8'd11;
        rom[107][3] = -8'd11;
        rom[107][4] = -8'd30;
        rom[107][5] = -8'd8;
        rom[107][6] = -8'd5;
        rom[107][7] = 8'd29;
        rom[107][8] = -8'd40;
        rom[107][9] = -8'd3;
        rom[107][10] = 8'd23;
        rom[107][11] = 8'd26;
        rom[107][12] = 8'd53;
        rom[107][13] = -8'd6;
        rom[107][14] = 8'd1;
        rom[107][15] = 8'd7;
        rom[107][16] = -8'd49;
        rom[107][17] = 8'd14;
        rom[107][18] = -8'd10;
        rom[107][19] = 8'd3;
        rom[107][20] = -8'd36;
        rom[107][21] = -8'd8;
        rom[107][22] = -8'd36;
        rom[107][23] = 8'd31;
        rom[107][24] = 8'd6;
        rom[107][25] = 8'd33;
        rom[107][26] = -8'd10;
        rom[107][27] = 8'd20;
        rom[107][28] = -8'd1;
        rom[107][29] = 8'd6;
        rom[107][30] = 8'd16;
        rom[107][31] = 8'd2;
        rom[108][0] = -8'd25;
        rom[108][1] = 8'd19;
        rom[108][2] = 8'd29;
        rom[108][3] = -8'd27;
        rom[108][4] = -8'd8;
        rom[108][5] = 8'd29;
        rom[108][6] = 8'd24;
        rom[108][7] = 8'd12;
        rom[108][8] = 8'd39;
        rom[108][9] = -8'd43;
        rom[108][10] = 8'd17;
        rom[108][11] = -8'd25;
        rom[108][12] = -8'd36;
        rom[108][13] = 8'd13;
        rom[108][14] = 8'd14;
        rom[108][15] = -8'd1;
        rom[108][16] = -8'd23;
        rom[108][17] = 8'd2;
        rom[108][18] = 8'd16;
        rom[108][19] = 8'd26;
        rom[108][20] = -8'd22;
        rom[108][21] = -8'd14;
        rom[108][22] = -8'd16;
        rom[108][23] = -8'd19;
        rom[108][24] = 8'd10;
        rom[108][25] = -8'd19;
        rom[108][26] = 8'd18;
        rom[108][27] = 8'd5;
        rom[108][28] = 8'd31;
        rom[108][29] = -8'd8;
        rom[108][30] = 8'd20;
        rom[108][31] = -8'd18;
        rom[109][0] = 8'd2;
        rom[109][1] = -8'd34;
        rom[109][2] = -8'd27;
        rom[109][3] = -8'd14;
        rom[109][4] = -8'd10;
        rom[109][5] = 8'd53;
        rom[109][6] = 8'd15;
        rom[109][7] = -8'd12;
        rom[109][8] = 8'd33;
        rom[109][9] = 8'd18;
        rom[109][10] = 8'd24;
        rom[109][11] = -8'd3;
        rom[109][12] = -8'd24;
        rom[109][13] = -8'd24;
        rom[109][14] = 8'd4;
        rom[109][15] = -8'd17;
        rom[109][16] = 8'd1;
        rom[109][17] = -8'd28;
        rom[109][18] = -8'd30;
        rom[109][19] = 8'd1;
        rom[109][20] = -8'd40;
        rom[109][21] = -8'd25;
        rom[109][22] = 8'd17;
        rom[109][23] = -8'd10;
        rom[109][24] = -8'd98;
        rom[109][25] = -8'd35;
        rom[109][26] = -8'd3;
        rom[109][27] = 8'd8;
        rom[109][28] = 8'd2;
        rom[109][29] = 8'd4;
        rom[109][30] = 8'd49;
        rom[109][31] = 8'd25;
        rom[110][0] = 8'd13;
        rom[110][1] = -8'd25;
        rom[110][2] = -8'd46;
        rom[110][3] = 8'd6;
        rom[110][4] = 8'd21;
        rom[110][5] = 8'd25;
        rom[110][6] = -8'd5;
        rom[110][7] = -8'd8;
        rom[110][8] = 8'd12;
        rom[110][9] = 8'd0;
        rom[110][10] = -8'd19;
        rom[110][11] = 8'd2;
        rom[110][12] = 8'd2;
        rom[110][13] = 8'd0;
        rom[110][14] = -8'd10;
        rom[110][15] = 8'd16;
        rom[110][16] = 8'd12;
        rom[110][17] = -8'd42;
        rom[110][18] = -8'd1;
        rom[110][19] = 8'd2;
        rom[110][20] = 8'd6;
        rom[110][21] = 8'd12;
        rom[110][22] = -8'd7;
        rom[110][23] = 8'd20;
        rom[110][24] = -8'd14;
        rom[110][25] = -8'd6;
        rom[110][26] = 8'd8;
        rom[110][27] = -8'd14;
        rom[110][28] = 8'd7;
        rom[110][29] = -8'd14;
        rom[110][30] = 8'd28;
        rom[110][31] = 8'd19;
        rom[111][0] = -8'd35;
        rom[111][1] = 8'd19;
        rom[111][2] = 8'd13;
        rom[111][3] = 8'd2;
        rom[111][4] = 8'd44;
        rom[111][5] = -8'd31;
        rom[111][6] = 8'd2;
        rom[111][7] = -8'd12;
        rom[111][8] = 8'd0;
        rom[111][9] = -8'd43;
        rom[111][10] = -8'd30;
        rom[111][11] = -8'd3;
        rom[111][12] = -8'd38;
        rom[111][13] = -8'd1;
        rom[111][14] = -8'd26;
        rom[111][15] = -8'd13;
        rom[111][16] = 8'd47;
        rom[111][17] = 8'd50;
        rom[111][18] = -8'd37;
        rom[111][19] = 8'd11;
        rom[111][20] = -8'd15;
        rom[111][21] = 8'd23;
        rom[111][22] = 8'd12;
        rom[111][23] = -8'd16;
        rom[111][24] = -8'd5;
        rom[111][25] = -8'd6;
        rom[111][26] = 8'd8;
        rom[111][27] = 8'd7;
        rom[111][28] = -8'd12;
        rom[111][29] = 8'd1;
        rom[111][30] = -8'd1;
        rom[111][31] = 8'd2;
        rom[112][0] = -8'd12;
        rom[112][1] = 8'd2;
        rom[112][2] = 8'd24;
        rom[112][3] = 8'd15;
        rom[112][4] = 8'd1;
        rom[112][5] = -8'd2;
        rom[112][6] = -8'd7;
        rom[112][7] = -8'd8;
        rom[112][8] = -8'd15;
        rom[112][9] = -8'd24;
        rom[112][10] = 8'd28;
        rom[112][11] = -8'd18;
        rom[112][12] = 8'd22;
        rom[112][13] = 8'd10;
        rom[112][14] = 8'd8;
        rom[112][15] = -8'd33;
        rom[112][16] = -8'd27;
        rom[112][17] = -8'd19;
        rom[112][18] = 8'd1;
        rom[112][19] = -8'd58;
        rom[112][20] = 8'd20;
        rom[112][21] = -8'd55;
        rom[112][22] = -8'd8;
        rom[112][23] = -8'd30;
        rom[112][24] = 8'd10;
        rom[112][25] = -8'd38;
        rom[112][26] = -8'd20;
        rom[112][27] = -8'd20;
        rom[112][28] = -8'd17;
        rom[112][29] = -8'd10;
        rom[112][30] = -8'd32;
        rom[112][31] = -8'd6;
        rom[113][0] = 8'd2;
        rom[113][1] = 8'd12;
        rom[113][2] = 8'd36;
        rom[113][3] = -8'd29;
        rom[113][4] = 8'd12;
        rom[113][5] = 8'd15;
        rom[113][6] = -8'd12;
        rom[113][7] = 8'd23;
        rom[113][8] = 8'd40;
        rom[113][9] = -8'd4;
        rom[113][10] = 8'd23;
        rom[113][11] = 8'd2;
        rom[113][12] = -8'd5;
        rom[113][13] = -8'd14;
        rom[113][14] = 8'd25;
        rom[113][15] = 8'd4;
        rom[113][16] = 8'd15;
        rom[113][17] = 8'd44;
        rom[113][18] = -8'd48;
        rom[113][19] = 8'd4;
        rom[113][20] = 8'd4;
        rom[113][21] = -8'd13;
        rom[113][22] = 8'd19;
        rom[113][23] = -8'd19;
        rom[113][24] = -8'd66;
        rom[113][25] = 8'd27;
        rom[113][26] = 8'd0;
        rom[113][27] = -8'd24;
        rom[113][28] = 8'd7;
        rom[113][29] = -8'd19;
        rom[113][30] = 8'd12;
        rom[113][31] = 8'd17;
        rom[114][0] = -8'd38;
        rom[114][1] = 8'd14;
        rom[114][2] = 8'd29;
        rom[114][3] = 8'd41;
        rom[114][4] = -8'd15;
        rom[114][5] = -8'd10;
        rom[114][6] = 8'd48;
        rom[114][7] = -8'd32;
        rom[114][8] = 8'd11;
        rom[114][9] = -8'd35;
        rom[114][10] = -8'd25;
        rom[114][11] = -8'd18;
        rom[114][12] = -8'd4;
        rom[114][13] = -8'd21;
        rom[114][14] = -8'd24;
        rom[114][15] = 8'd22;
        rom[114][16] = 8'd49;
        rom[114][17] = -8'd11;
        rom[114][18] = 8'd27;
        rom[114][19] = -8'd3;
        rom[114][20] = -8'd24;
        rom[114][21] = 8'd19;
        rom[114][22] = 8'd20;
        rom[114][23] = -8'd31;
        rom[114][24] = -8'd11;
        rom[114][25] = -8'd11;
        rom[114][26] = -8'd16;
        rom[114][27] = 8'd5;
        rom[114][28] = 8'd35;
        rom[114][29] = 8'd8;
        rom[114][30] = -8'd11;
        rom[114][31] = 8'd5;
        rom[115][0] = 8'd5;
        rom[115][1] = -8'd38;
        rom[115][2] = -8'd66;
        rom[115][3] = 8'd24;
        rom[115][4] = -8'd10;
        rom[115][5] = 8'd29;
        rom[115][6] = 8'd6;
        rom[115][7] = 8'd1;
        rom[115][8] = 8'd22;
        rom[115][9] = 8'd0;
        rom[115][10] = -8'd25;
        rom[115][11] = -8'd13;
        rom[115][12] = 8'd9;
        rom[115][13] = 8'd36;
        rom[115][14] = 8'd20;
        rom[115][15] = 8'd12;
        rom[115][16] = -8'd4;
        rom[115][17] = -8'd24;
        rom[115][18] = 8'd14;
        rom[115][19] = -8'd3;
        rom[115][20] = 8'd6;
        rom[115][21] = 8'd6;
        rom[115][22] = 8'd14;
        rom[115][23] = -8'd5;
        rom[115][24] = -8'd26;
        rom[115][25] = -8'd24;
        rom[115][26] = 8'd10;
        rom[115][27] = -8'd20;
        rom[115][28] = -8'd2;
        rom[115][29] = -8'd14;
        rom[115][30] = -8'd2;
        rom[115][31] = -8'd44;
        rom[116][0] = 8'd51;
        rom[116][1] = 8'd8;
        rom[116][2] = 8'd21;
        rom[116][3] = -8'd11;
        rom[116][4] = 8'd47;
        rom[116][5] = -8'd24;
        rom[116][6] = -8'd6;
        rom[116][7] = -8'd8;
        rom[116][8] = -8'd38;
        rom[116][9] = 8'd11;
        rom[116][10] = 8'd25;
        rom[116][11] = 8'd14;
        rom[116][12] = 8'd26;
        rom[116][13] = -8'd10;
        rom[116][14] = 8'd4;
        rom[116][15] = -8'd25;
        rom[116][16] = 8'd5;
        rom[116][17] = 8'd6;
        rom[116][18] = -8'd8;
        rom[116][19] = -8'd41;
        rom[116][20] = -8'd9;
        rom[116][21] = 8'd19;
        rom[116][22] = -8'd65;
        rom[116][23] = 8'd18;
        rom[116][24] = 8'd11;
        rom[116][25] = 8'd10;
        rom[116][26] = -8'd28;
        rom[116][27] = 8'd27;
        rom[116][28] = -8'd1;
        rom[116][29] = -8'd18;
        rom[116][30] = -8'd41;
        rom[116][31] = -8'd24;
        rom[117][0] = -8'd7;
        rom[117][1] = 8'd9;
        rom[117][2] = 8'd3;
        rom[117][3] = 8'd2;
        rom[117][4] = -8'd3;
        rom[117][5] = 8'd31;
        rom[117][6] = 8'd1;
        rom[117][7] = 8'd3;
        rom[117][8] = 8'd41;
        rom[117][9] = -8'd9;
        rom[117][10] = -8'd20;
        rom[117][11] = -8'd44;
        rom[117][12] = -8'd22;
        rom[117][13] = 8'd7;
        rom[117][14] = -8'd16;
        rom[117][15] = -8'd26;
        rom[117][16] = -8'd36;
        rom[117][17] = -8'd21;
        rom[117][18] = -8'd16;
        rom[117][19] = 8'd5;
        rom[117][20] = 8'd14;
        rom[117][21] = 8'd11;
        rom[117][22] = 8'd13;
        rom[117][23] = -8'd5;
        rom[117][24] = 8'd15;
        rom[117][25] = 8'd2;
        rom[117][26] = -8'd26;
        rom[117][27] = 8'd7;
        rom[117][28] = 8'd1;
        rom[117][29] = 8'd4;
        rom[117][30] = 8'd12;
        rom[117][31] = -8'd8;
        rom[118][0] = -8'd23;
        rom[118][1] = -8'd15;
        rom[118][2] = -8'd23;
        rom[118][3] = 8'd26;
        rom[118][4] = 8'd2;
        rom[118][5] = 8'd13;
        rom[118][6] = -8'd19;
        rom[118][7] = 8'd8;
        rom[118][8] = 8'd30;
        rom[118][9] = 8'd25;
        rom[118][10] = 8'd12;
        rom[118][11] = 8'd3;
        rom[118][12] = 8'd3;
        rom[118][13] = 8'd4;
        rom[118][14] = 8'd22;
        rom[118][15] = 8'd3;
        rom[118][16] = 8'd2;
        rom[118][17] = 8'd42;
        rom[118][18] = -8'd17;
        rom[118][19] = 8'd17;
        rom[118][20] = -8'd12;
        rom[118][21] = -8'd25;
        rom[118][22] = -8'd6;
        rom[118][23] = 8'd0;
        rom[118][24] = -8'd34;
        rom[118][25] = -8'd2;
        rom[118][26] = -8'd15;
        rom[118][27] = -8'd31;
        rom[118][28] = -8'd10;
        rom[118][29] = 8'd0;
        rom[118][30] = -8'd1;
        rom[118][31] = 8'd12;
        rom[119][0] = 8'd8;
        rom[119][1] = -8'd34;
        rom[119][2] = 8'd12;
        rom[119][3] = 8'd6;
        rom[119][4] = 8'd12;
        rom[119][5] = 8'd31;
        rom[119][6] = -8'd15;
        rom[119][7] = 8'd4;
        rom[119][8] = -8'd47;
        rom[119][9] = 8'd17;
        rom[119][10] = -8'd32;
        rom[119][11] = 8'd8;
        rom[119][12] = -8'd6;
        rom[119][13] = -8'd14;
        rom[119][14] = 8'd38;
        rom[119][15] = -8'd21;
        rom[119][16] = 8'd18;
        rom[119][17] = 8'd32;
        rom[119][18] = -8'd29;
        rom[119][19] = 8'd3;
        rom[119][20] = 8'd8;
        rom[119][21] = -8'd17;
        rom[119][22] = -8'd30;
        rom[119][23] = 8'd26;
        rom[119][24] = -8'd8;
        rom[119][25] = 8'd4;
        rom[119][26] = -8'd5;
        rom[119][27] = -8'd4;
        rom[119][28] = 8'd24;
        rom[119][29] = -8'd1;
        rom[119][30] = -8'd4;
        rom[119][31] = 8'd7;
        rom[120][0] = -8'd36;
        rom[120][1] = -8'd6;
        rom[120][2] = -8'd7;
        rom[120][3] = -8'd25;
        rom[120][4] = -8'd61;
        rom[120][5] = 8'd0;
        rom[120][6] = -8'd7;
        rom[120][7] = -8'd14;
        rom[120][8] = -8'd5;
        rom[120][9] = -8'd18;
        rom[120][10] = -8'd30;
        rom[120][11] = -8'd51;
        rom[120][12] = -8'd17;
        rom[120][13] = 8'd43;
        rom[120][14] = 8'd3;
        rom[120][15] = -8'd17;
        rom[120][16] = -8'd30;
        rom[120][17] = -8'd58;
        rom[120][18] = 8'd23;
        rom[120][19] = -8'd30;
        rom[120][20] = 8'd58;
        rom[120][21] = 8'd45;
        rom[120][22] = -8'd32;
        rom[120][23] = -8'd20;
        rom[120][24] = 8'd10;
        rom[120][25] = -8'd10;
        rom[120][26] = -8'd18;
        rom[120][27] = -8'd2;
        rom[120][28] = -8'd1;
        rom[120][29] = 8'd4;
        rom[120][30] = -8'd63;
        rom[120][31] = 8'd2;
        rom[121][0] = -8'd19;
        rom[121][1] = 8'd14;
        rom[121][2] = -8'd29;
        rom[121][3] = -8'd2;
        rom[121][4] = -8'd20;
        rom[121][5] = 8'd62;
        rom[121][6] = 8'd40;
        rom[121][7] = 8'd39;
        rom[121][8] = 8'd2;
        rom[121][9] = 8'd7;
        rom[121][10] = 8'd0;
        rom[121][11] = -8'd16;
        rom[121][12] = -8'd12;
        rom[121][13] = 8'd15;
        rom[121][14] = 8'd11;
        rom[121][15] = 8'd18;
        rom[121][16] = 8'd13;
        rom[121][17] = 8'd19;
        rom[121][18] = -8'd24;
        rom[121][19] = 8'd10;
        rom[121][20] = 8'd6;
        rom[121][21] = 8'd9;
        rom[121][22] = 8'd11;
        rom[121][23] = -8'd7;
        rom[121][24] = 8'd19;
        rom[121][25] = -8'd47;
        rom[121][26] = -8'd1;
        rom[121][27] = 8'd12;
        rom[121][28] = 8'd23;
        rom[121][29] = -8'd1;
        rom[121][30] = -8'd57;
        rom[121][31] = 8'd30;
        rom[122][0] = -8'd21;
        rom[122][1] = -8'd8;
        rom[122][2] = 8'd20;
        rom[122][3] = 8'd0;
        rom[122][4] = 8'd5;
        rom[122][5] = 8'd38;
        rom[122][6] = -8'd19;
        rom[122][7] = -8'd6;
        rom[122][8] = 8'd0;
        rom[122][9] = 8'd0;
        rom[122][10] = -8'd17;
        rom[122][11] = -8'd31;
        rom[122][12] = -8'd23;
        rom[122][13] = -8'd30;
        rom[122][14] = -8'd24;
        rom[122][15] = 8'd12;
        rom[122][16] = 8'd3;
        rom[122][17] = -8'd12;
        rom[122][18] = -8'd10;
        rom[122][19] = 8'd12;
        rom[122][20] = 8'd17;
        rom[122][21] = -8'd3;
        rom[122][22] = 8'd2;
        rom[122][23] = 8'd23;
        rom[122][24] = 8'd10;
        rom[122][25] = -8'd32;
        rom[122][26] = 8'd0;
        rom[122][27] = -8'd11;
        rom[122][28] = -8'd10;
        rom[122][29] = 8'd2;
        rom[122][30] = 8'd3;
        rom[122][31] = 8'd7;
        rom[123][0] = 8'd0;
        rom[123][1] = 8'd2;
        rom[123][2] = -8'd20;
        rom[123][3] = -8'd6;
        rom[123][4] = 8'd8;
        rom[123][5] = 8'd6;
        rom[123][6] = -8'd9;
        rom[123][7] = 8'd26;
        rom[123][8] = -8'd10;
        rom[123][9] = -8'd12;
        rom[123][10] = 8'd14;
        rom[123][11] = 8'd43;
        rom[123][12] = 8'd21;
        rom[123][13] = 8'd10;
        rom[123][14] = -8'd45;
        rom[123][15] = -8'd7;
        rom[123][16] = -8'd10;
        rom[123][17] = -8'd41;
        rom[123][18] = 8'd24;
        rom[123][19] = -8'd14;
        rom[123][20] = 8'd4;
        rom[123][21] = 8'd27;
        rom[123][22] = -8'd12;
        rom[123][23] = 8'd27;
        rom[123][24] = -8'd30;
        rom[123][25] = -8'd14;
        rom[123][26] = 8'd13;
        rom[123][27] = -8'd38;
        rom[123][28] = 8'd12;
        rom[123][29] = -8'd13;
        rom[123][30] = 8'd17;
        rom[123][31] = 8'd21;
        rom[124][0] = -8'd4;
        rom[124][1] = 8'd5;
        rom[124][2] = 8'd11;
        rom[124][3] = -8'd16;
        rom[124][4] = 8'd3;
        rom[124][5] = 8'd4;
        rom[124][6] = 8'd30;
        rom[124][7] = 8'd26;
        rom[124][8] = 8'd29;
        rom[124][9] = -8'd16;
        rom[124][10] = -8'd3;
        rom[124][11] = 8'd16;
        rom[124][12] = -8'd33;
        rom[124][13] = -8'd40;
        rom[124][14] = 8'd20;
        rom[124][15] = -8'd19;
        rom[124][16] = -8'd32;
        rom[124][17] = 8'd4;
        rom[124][18] = 8'd29;
        rom[124][19] = 8'd3;
        rom[124][20] = -8'd52;
        rom[124][21] = -8'd4;
        rom[124][22] = -8'd16;
        rom[124][23] = -8'd80;
        rom[124][24] = -8'd12;
        rom[124][25] = -8'd17;
        rom[124][26] = -8'd11;
        rom[124][27] = 8'd52;
        rom[124][28] = -8'd9;
        rom[124][29] = 8'd7;
        rom[124][30] = -8'd17;
        rom[124][31] = -8'd29;
        rom[125][0] = 8'd14;
        rom[125][1] = -8'd10;
        rom[125][2] = 8'd15;
        rom[125][3] = 8'd2;
        rom[125][4] = 8'd30;
        rom[125][5] = 8'd3;
        rom[125][6] = 8'd40;
        rom[125][7] = -8'd70;
        rom[125][8] = -8'd2;
        rom[125][9] = 8'd43;
        rom[125][10] = 8'd1;
        rom[125][11] = -8'd30;
        rom[125][12] = 8'd21;
        rom[125][13] = -8'd8;
        rom[125][14] = -8'd45;
        rom[125][15] = 8'd21;
        rom[125][16] = 8'd40;
        rom[125][17] = -8'd12;
        rom[125][18] = 8'd2;
        rom[125][19] = 8'd29;
        rom[125][20] = 8'd17;
        rom[125][21] = 8'd2;
        rom[125][22] = -8'd25;
        rom[125][23] = 8'd0;
        rom[125][24] = -8'd33;
        rom[125][25] = 8'd30;
        rom[125][26] = -8'd4;
        rom[125][27] = -8'd7;
        rom[125][28] = -8'd5;
        rom[125][29] = 8'd0;
        rom[125][30] = -8'd1;
        rom[125][31] = -8'd18;
        rom[126][0] = 8'd22;
        rom[126][1] = 8'd11;
        rom[126][2] = -8'd1;
        rom[126][3] = -8'd13;
        rom[126][4] = -8'd28;
        rom[126][5] = 8'd17;
        rom[126][6] = 8'd8;
        rom[126][7] = -8'd5;
        rom[126][8] = 8'd11;
        rom[126][9] = -8'd34;
        rom[126][10] = -8'd6;
        rom[126][11] = 8'd37;
        rom[126][12] = -8'd5;
        rom[126][13] = -8'd19;
        rom[126][14] = 8'd17;
        rom[126][15] = 8'd29;
        rom[126][16] = -8'd12;
        rom[126][17] = 8'd13;
        rom[126][18] = 8'd32;
        rom[126][19] = 8'd4;
        rom[126][20] = -8'd13;
        rom[126][21] = 8'd33;
        rom[126][22] = -8'd60;
        rom[126][23] = -8'd47;
        rom[126][24] = 8'd29;
        rom[126][25] = 8'd31;
        rom[126][26] = 8'd4;
        rom[126][27] = -8'd8;
        rom[126][28] = 8'd25;
        rom[126][29] = -8'd12;
        rom[126][30] = -8'd19;
        rom[126][31] = -8'd29;
        rom[127][0] = -8'd40;
        rom[127][1] = 8'd10;
        rom[127][2] = 8'd42;
        rom[127][3] = 8'd1;
        rom[127][4] = 8'd30;
        rom[127][5] = 8'd16;
        rom[127][6] = -8'd9;
        rom[127][7] = 8'd17;
        rom[127][8] = -8'd1;
        rom[127][9] = -8'd61;
        rom[127][10] = -8'd25;
        rom[127][11] = -8'd22;
        rom[127][12] = 8'd38;
        rom[127][13] = 8'd14;
        rom[127][14] = -8'd58;
        rom[127][15] = 8'd22;
        rom[127][16] = -8'd9;
        rom[127][17] = 8'd17;
        rom[127][18] = 8'd10;
        rom[127][19] = -8'd20;
        rom[127][20] = -8'd39;
        rom[127][21] = 8'd35;
        rom[127][22] = -8'd2;
        rom[127][23] = -8'd11;
        rom[127][24] = -8'd30;
        rom[127][25] = -8'd15;
        rom[127][26] = -8'd21;
        rom[127][27] = 8'd1;
        rom[127][28] = -8'd59;
        rom[127][29] = 8'd7;
        rom[127][30] = 8'd6;
        rom[127][31] = -8'd40;
        rom[128][0] = -8'd6;
        rom[128][1] = 8'd22;
        rom[128][2] = -8'd12;
        rom[128][3] = -8'd39;
        rom[128][4] = 8'd20;
        rom[128][5] = 8'd0;
        rom[128][6] = 8'd6;
        rom[128][7] = -8'd26;
        rom[128][8] = 8'd22;
        rom[128][9] = -8'd23;
        rom[128][10] = 8'd23;
        rom[128][11] = 8'd13;
        rom[128][12] = -8'd12;
        rom[128][13] = 8'd9;
        rom[128][14] = 8'd5;
        rom[128][15] = -8'd63;
        rom[128][16] = -8'd29;
        rom[128][17] = 8'd13;
        rom[128][18] = -8'd18;
        rom[128][19] = -8'd19;
        rom[128][20] = -8'd49;
        rom[128][21] = -8'd34;
        rom[128][22] = 8'd9;
        rom[128][23] = 8'd7;
        rom[128][24] = 8'd1;
        rom[128][25] = 8'd19;
        rom[128][26] = -8'd4;
        rom[128][27] = 8'd3;
        rom[128][28] = -8'd6;
        rom[128][29] = -8'd9;
        rom[128][30] = 8'd23;
        rom[128][31] = 8'd23;
        rom[129][0] = 8'd15;
        rom[129][1] = -8'd28;
        rom[129][2] = -8'd23;
        rom[129][3] = -8'd44;
        rom[129][4] = -8'd81;
        rom[129][5] = 8'd22;
        rom[129][6] = -8'd29;
        rom[129][7] = 8'd3;
        rom[129][8] = -8'd43;
        rom[129][9] = -8'd6;
        rom[129][10] = -8'd11;
        rom[129][11] = -8'd9;
        rom[129][12] = -8'd18;
        rom[129][13] = -8'd13;
        rom[129][14] = 8'd3;
        rom[129][15] = 8'd0;
        rom[129][16] = 8'd53;
        rom[129][17] = -8'd18;
        rom[129][18] = 8'd14;
        rom[129][19] = -8'd6;
        rom[129][20] = 8'd13;
        rom[129][21] = 8'd28;
        rom[129][22] = -8'd28;
        rom[129][23] = -8'd14;
        rom[129][24] = 8'd28;
        rom[129][25] = -8'd28;
        rom[129][26] = -8'd5;
        rom[129][27] = 8'd20;
        rom[129][28] = 8'd6;
        rom[129][29] = -8'd12;
        rom[129][30] = -8'd62;
        rom[129][31] = -8'd44;
        rom[130][0] = -8'd38;
        rom[130][1] = -8'd20;
        rom[130][2] = -8'd29;
        rom[130][3] = 8'd10;
        rom[130][4] = -8'd4;
        rom[130][5] = 8'd27;
        rom[130][6] = 8'd14;
        rom[130][7] = 8'd0;
        rom[130][8] = -8'd20;
        rom[130][9] = -8'd32;
        rom[130][10] = -8'd25;
        rom[130][11] = -8'd43;
        rom[130][12] = -8'd20;
        rom[130][13] = -8'd53;
        rom[130][14] = -8'd18;
        rom[130][15] = -8'd32;
        rom[130][16] = -8'd45;
        rom[130][17] = 8'd22;
        rom[130][18] = -8'd9;
        rom[130][19] = -8'd68;
        rom[130][20] = -8'd20;
        rom[130][21] = -8'd31;
        rom[130][22] = 8'd45;
        rom[130][23] = 8'd10;
        rom[130][24] = -8'd3;
        rom[130][25] = -8'd57;
        rom[130][26] = -8'd23;
        rom[130][27] = -8'd89;
        rom[130][28] = -8'd28;
        rom[130][29] = -8'd1;
        rom[130][30] = 8'd3;
        rom[130][31] = -8'd5;
        rom[131][0] = 8'd6;
        rom[131][1] = -8'd25;
        rom[131][2] = 8'd18;
        rom[131][3] = 8'd16;
        rom[131][4] = -8'd35;
        rom[131][5] = -8'd11;
        rom[131][6] = 8'd28;
        rom[131][7] = -8'd5;
        rom[131][8] = -8'd30;
        rom[131][9] = -8'd41;
        rom[131][10] = -8'd30;
        rom[131][11] = 8'd27;
        rom[131][12] = 8'd2;
        rom[131][13] = -8'd28;
        rom[131][14] = 8'd3;
        rom[131][15] = -8'd46;
        rom[131][16] = -8'd13;
        rom[131][17] = -8'd3;
        rom[131][18] = -8'd7;
        rom[131][19] = 8'd18;
        rom[131][20] = 8'd24;
        rom[131][21] = -8'd38;
        rom[131][22] = 8'd25;
        rom[131][23] = -8'd9;
        rom[131][24] = 8'd45;
        rom[131][25] = 8'd31;
        rom[131][26] = 8'd3;
        rom[131][27] = 8'd0;
        rom[131][28] = -8'd58;
        rom[131][29] = -8'd12;
        rom[131][30] = 8'd24;
        rom[131][31] = -8'd24;
        rom[132][0] = -8'd2;
        rom[132][1] = -8'd41;
        rom[132][2] = 8'd34;
        rom[132][3] = 8'd15;
        rom[132][4] = 8'd5;
        rom[132][5] = 8'd27;
        rom[132][6] = 8'd4;
        rom[132][7] = 8'd39;
        rom[132][8] = -8'd7;
        rom[132][9] = -8'd36;
        rom[132][10] = 8'd19;
        rom[132][11] = 8'd39;
        rom[132][12] = -8'd12;
        rom[132][13] = -8'd5;
        rom[132][14] = 8'd18;
        rom[132][15] = 8'd35;
        rom[132][16] = 8'd0;
        rom[132][17] = -8'd23;
        rom[132][18] = 8'd17;
        rom[132][19] = -8'd49;
        rom[132][20] = 8'd26;
        rom[132][21] = -8'd3;
        rom[132][22] = -8'd36;
        rom[132][23] = -8'd28;
        rom[132][24] = 8'd26;
        rom[132][25] = -8'd52;
        rom[132][26] = -8'd46;
        rom[132][27] = -8'd9;
        rom[132][28] = 8'd10;
        rom[132][29] = -8'd11;
        rom[132][30] = -8'd7;
        rom[132][31] = 8'd18;
        rom[133][0] = -8'd45;
        rom[133][1] = -8'd21;
        rom[133][2] = -8'd35;
        rom[133][3] = -8'd21;
        rom[133][4] = -8'd54;
        rom[133][5] = 8'd29;
        rom[133][6] = 8'd2;
        rom[133][7] = -8'd11;
        rom[133][8] = 8'd16;
        rom[133][9] = -8'd1;
        rom[133][10] = 8'd7;
        rom[133][11] = -8'd31;
        rom[133][12] = -8'd63;
        rom[133][13] = 8'd29;
        rom[133][14] = 8'd37;
        rom[133][15] = -8'd87;
        rom[133][16] = -8'd12;
        rom[133][17] = 8'd24;
        rom[133][18] = -8'd61;
        rom[133][19] = 8'd28;
        rom[133][20] = -8'd25;
        rom[133][21] = 8'd3;
        rom[133][22] = -8'd17;
        rom[133][23] = 8'd1;
        rom[133][24] = 8'd16;
        rom[133][25] = -8'd20;
        rom[133][26] = -8'd20;
        rom[133][27] = -8'd12;
        rom[133][28] = -8'd28;
        rom[133][29] = -8'd5;
        rom[133][30] = -8'd8;
        rom[133][31] = -8'd28;
        rom[134][0] = -8'd27;
        rom[134][1] = 8'd4;
        rom[134][2] = -8'd8;
        rom[134][3] = -8'd27;
        rom[134][4] = -8'd27;
        rom[134][5] = 8'd39;
        rom[134][6] = 8'd17;
        rom[134][7] = -8'd51;
        rom[134][8] = 8'd29;
        rom[134][9] = -8'd48;
        rom[134][10] = -8'd44;
        rom[134][11] = -8'd11;
        rom[134][12] = -8'd16;
        rom[134][13] = 8'd23;
        rom[134][14] = -8'd10;
        rom[134][15] = -8'd23;
        rom[134][16] = 8'd31;
        rom[134][17] = 8'd6;
        rom[134][18] = -8'd63;
        rom[134][19] = -8'd8;
        rom[134][20] = -8'd8;
        rom[134][21] = -8'd12;
        rom[134][22] = 8'd10;
        rom[134][23] = 8'd13;
        rom[134][24] = 8'd4;
        rom[134][25] = -8'd33;
        rom[134][26] = 8'd17;
        rom[134][27] = -8'd16;
        rom[134][28] = 8'd22;
        rom[134][29] = -8'd4;
        rom[134][30] = -8'd40;
        rom[134][31] = 8'd40;
        rom[135][0] = 8'd9;
        rom[135][1] = 8'd14;
        rom[135][2] = -8'd17;
        rom[135][3] = -8'd20;
        rom[135][4] = 8'd6;
        rom[135][5] = -8'd28;
        rom[135][6] = -8'd12;
        rom[135][7] = 8'd10;
        rom[135][8] = 8'd16;
        rom[135][9] = 8'd6;
        rom[135][10] = 8'd33;
        rom[135][11] = -8'd3;
        rom[135][12] = 8'd47;
        rom[135][13] = 8'd9;
        rom[135][14] = -8'd60;
        rom[135][15] = 8'd0;
        rom[135][16] = 8'd3;
        rom[135][17] = -8'd3;
        rom[135][18] = 8'd1;
        rom[135][19] = 8'd1;
        rom[135][20] = -8'd24;
        rom[135][21] = -8'd9;
        rom[135][22] = -8'd9;
        rom[135][23] = -8'd14;
        rom[135][24] = 8'd13;
        rom[135][25] = 8'd22;
        rom[135][26] = 8'd30;
        rom[135][27] = 8'd13;
        rom[135][28] = -8'd12;
        rom[135][29] = -8'd7;
        rom[135][30] = -8'd20;
        rom[135][31] = 8'd12;
        rom[136][0] = -8'd11;
        rom[136][1] = 8'd26;
        rom[136][2] = 8'd11;
        rom[136][3] = 8'd11;
        rom[136][4] = -8'd18;
        rom[136][5] = 8'd8;
        rom[136][6] = 8'd31;
        rom[136][7] = 8'd7;
        rom[136][8] = -8'd17;
        rom[136][9] = 8'd4;
        rom[136][10] = -8'd7;
        rom[136][11] = 8'd28;
        rom[136][12] = -8'd22;
        rom[136][13] = -8'd7;
        rom[136][14] = -8'd9;
        rom[136][15] = -8'd26;
        rom[136][16] = -8'd30;
        rom[136][17] = -8'd28;
        rom[136][18] = -8'd2;
        rom[136][19] = -8'd44;
        rom[136][20] = 8'd5;
        rom[136][21] = 8'd8;
        rom[136][22] = 8'd6;
        rom[136][23] = 8'd1;
        rom[136][24] = 8'd26;
        rom[136][25] = 8'd0;
        rom[136][26] = -8'd6;
        rom[136][27] = 8'd3;
        rom[136][28] = -8'd29;
        rom[136][29] = 8'd1;
        rom[136][30] = -8'd16;
        rom[136][31] = 8'd8;
        rom[137][0] = -8'd3;
        rom[137][1] = -8'd11;
        rom[137][2] = -8'd4;
        rom[137][3] = -8'd19;
        rom[137][4] = -8'd5;
        rom[137][5] = 8'd36;
        rom[137][6] = -8'd5;
        rom[137][7] = -8'd40;
        rom[137][8] = -8'd35;
        rom[137][9] = -8'd9;
        rom[137][10] = 8'd3;
        rom[137][11] = -8'd26;
        rom[137][12] = 8'd19;
        rom[137][13] = -8'd24;
        rom[137][14] = -8'd32;
        rom[137][15] = 8'd22;
        rom[137][16] = -8'd40;
        rom[137][17] = -8'd1;
        rom[137][18] = -8'd13;
        rom[137][19] = -8'd38;
        rom[137][20] = -8'd25;
        rom[137][21] = -8'd34;
        rom[137][22] = 8'd7;
        rom[137][23] = 8'd38;
        rom[137][24] = 8'd16;
        rom[137][25] = 8'd0;
        rom[137][26] = -8'd17;
        rom[137][27] = -8'd54;
        rom[137][28] = -8'd18;
        rom[137][29] = 8'd6;
        rom[137][30] = 8'd8;
        rom[137][31] = -8'd4;
        rom[138][0] = -8'd22;
        rom[138][1] = -8'd35;
        rom[138][2] = -8'd17;
        rom[138][3] = -8'd37;
        rom[138][4] = -8'd18;
        rom[138][5] = -8'd38;
        rom[138][6] = -8'd11;
        rom[138][7] = 8'd13;
        rom[138][8] = 8'd19;
        rom[138][9] = -8'd5;
        rom[138][10] = -8'd22;
        rom[138][11] = 8'd48;
        rom[138][12] = -8'd41;
        rom[138][13] = -8'd54;
        rom[138][14] = 8'd1;
        rom[138][15] = 8'd32;
        rom[138][16] = 8'd18;
        rom[138][17] = 8'd53;
        rom[138][18] = 8'd16;
        rom[138][19] = -8'd24;
        rom[138][20] = -8'd10;
        rom[138][21] = 8'd26;
        rom[138][22] = -8'd8;
        rom[138][23] = 8'd17;
        rom[138][24] = 8'd10;
        rom[138][25] = -8'd38;
        rom[138][26] = 8'd9;
        rom[138][27] = -8'd84;
        rom[138][28] = -8'd17;
        rom[138][29] = -8'd10;
        rom[138][30] = 8'd17;
        rom[138][31] = -8'd50;
        rom[139][0] = 8'd21;
        rom[139][1] = 8'd1;
        rom[139][2] = -8'd17;
        rom[139][3] = -8'd20;
        rom[139][4] = -8'd45;
        rom[139][5] = -8'd2;
        rom[139][6] = -8'd42;
        rom[139][7] = 8'd1;
        rom[139][8] = 8'd2;
        rom[139][9] = 8'd33;
        rom[139][10] = -8'd8;
        rom[139][11] = -8'd23;
        rom[139][12] = -8'd4;
        rom[139][13] = 8'd5;
        rom[139][14] = 8'd11;
        rom[139][15] = 8'd24;
        rom[139][16] = -8'd10;
        rom[139][17] = 8'd3;
        rom[139][18] = 8'd16;
        rom[139][19] = 8'd7;
        rom[139][20] = 8'd23;
        rom[139][21] = 8'd31;
        rom[139][22] = -8'd25;
        rom[139][23] = 8'd45;
        rom[139][24] = 8'd32;
        rom[139][25] = 8'd17;
        rom[139][26] = 8'd16;
        rom[139][27] = 8'd3;
        rom[139][28] = 8'd11;
        rom[139][29] = -8'd10;
        rom[139][30] = -8'd33;
        rom[139][31] = -8'd26;
        rom[140][0] = 8'd3;
        rom[140][1] = -8'd21;
        rom[140][2] = -8'd7;
        rom[140][3] = -8'd30;
        rom[140][4] = -8'd38;
        rom[140][5] = 8'd13;
        rom[140][6] = 8'd12;
        rom[140][7] = -8'd45;
        rom[140][8] = -8'd23;
        rom[140][9] = -8'd42;
        rom[140][10] = 8'd24;
        rom[140][11] = 8'd5;
        rom[140][12] = -8'd17;
        rom[140][13] = -8'd17;
        rom[140][14] = 8'd2;
        rom[140][15] = -8'd13;
        rom[140][16] = -8'd4;
        rom[140][17] = 8'd6;
        rom[140][18] = 8'd12;
        rom[140][19] = 8'd15;
        rom[140][20] = -8'd47;
        rom[140][21] = -8'd39;
        rom[140][22] = 8'd7;
        rom[140][23] = 8'd23;
        rom[140][24] = 8'd36;
        rom[140][25] = 8'd5;
        rom[140][26] = 8'd3;
        rom[140][27] = 8'd5;
        rom[140][28] = -8'd53;
        rom[140][29] = -8'd3;
        rom[140][30] = -8'd7;
        rom[140][31] = -8'd45;
        rom[141][0] = 8'd30;
        rom[141][1] = -8'd51;
        rom[141][2] = -8'd14;
        rom[141][3] = -8'd6;
        rom[141][4] = 8'd0;
        rom[141][5] = 8'd61;
        rom[141][6] = -8'd60;
        rom[141][7] = -8'd6;
        rom[141][8] = -8'd12;
        rom[141][9] = 8'd8;
        rom[141][10] = 8'd22;
        rom[141][11] = 8'd12;
        rom[141][12] = -8'd19;
        rom[141][13] = -8'd28;
        rom[141][14] = 8'd2;
        rom[141][15] = -8'd20;
        rom[141][16] = -8'd40;
        rom[141][17] = -8'd42;
        rom[141][18] = -8'd53;
        rom[141][19] = -8'd10;
        rom[141][20] = -8'd43;
        rom[141][21] = -8'd7;
        rom[141][22] = 8'd20;
        rom[141][23] = -8'd1;
        rom[141][24] = 8'd9;
        rom[141][25] = 8'd18;
        rom[141][26] = 8'd11;
        rom[141][27] = -8'd9;
        rom[141][28] = -8'd19;
        rom[141][29] = -8'd7;
        rom[141][30] = 8'd30;
        rom[141][31] = -8'd6;
        rom[142][0] = 8'd35;
        rom[142][1] = -8'd1;
        rom[142][2] = -8'd21;
        rom[142][3] = -8'd19;
        rom[142][4] = 8'd21;
        rom[142][5] = 8'd34;
        rom[142][6] = -8'd28;
        rom[142][7] = -8'd13;
        rom[142][8] = -8'd2;
        rom[142][9] = 8'd6;
        rom[142][10] = 8'd11;
        rom[142][11] = -8'd13;
        rom[142][12] = 8'd3;
        rom[142][13] = 8'd11;
        rom[142][14] = -8'd35;
        rom[142][15] = 8'd30;
        rom[142][16] = -8'd20;
        rom[142][17] = -8'd50;
        rom[142][18] = -8'd10;
        rom[142][19] = 8'd4;
        rom[142][20] = -8'd16;
        rom[142][21] = -8'd9;
        rom[142][22] = -8'd16;
        rom[142][23] = -8'd37;
        rom[142][24] = -8'd18;
        rom[142][25] = 8'd19;
        rom[142][26] = -8'd6;
        rom[142][27] = 8'd1;
        rom[142][28] = -8'd1;
        rom[142][29] = -8'd12;
        rom[142][30] = 8'd20;
        rom[142][31] = 8'd26;
        rom[143][0] = 8'd4;
        rom[143][1] = 8'd9;
        rom[143][2] = -8'd5;
        rom[143][3] = -8'd22;
        rom[143][4] = -8'd1;
        rom[143][5] = 8'd6;
        rom[143][6] = 8'd2;
        rom[143][7] = -8'd10;
        rom[143][8] = 8'd1;
        rom[143][9] = -8'd78;
        rom[143][10] = -8'd33;
        rom[143][11] = 8'd39;
        rom[143][12] = -8'd22;
        rom[143][13] = -8'd19;
        rom[143][14] = -8'd44;
        rom[143][15] = -8'd40;
        rom[143][16] = -8'd2;
        rom[143][17] = 8'd1;
        rom[143][18] = -8'd22;
        rom[143][19] = -8'd4;
        rom[143][20] = -8'd62;
        rom[143][21] = -8'd31;
        rom[143][22] = 8'd16;
        rom[143][23] = -8'd16;
        rom[143][24] = -8'd8;
        rom[143][25] = -8'd21;
        rom[143][26] = -8'd20;
        rom[143][27] = -8'd18;
        rom[143][28] = -8'd66;
        rom[143][29] = -8'd5;
        rom[143][30] = 8'd15;
        rom[143][31] = 8'd14;
        rom[144][0] = -8'd17;
        rom[144][1] = 8'd1;
        rom[144][2] = 8'd18;
        rom[144][3] = -8'd4;
        rom[144][4] = -8'd26;
        rom[144][5] = 8'd8;
        rom[144][6] = 8'd16;
        rom[144][7] = 8'd1;
        rom[144][8] = -8'd2;
        rom[144][9] = 8'd1;
        rom[144][10] = 8'd29;
        rom[144][11] = -8'd5;
        rom[144][12] = 8'd36;
        rom[144][13] = -8'd14;
        rom[144][14] = 8'd15;
        rom[144][15] = -8'd27;
        rom[144][16] = -8'd26;
        rom[144][17] = -8'd2;
        rom[144][18] = 8'd11;
        rom[144][19] = -8'd103;
        rom[144][20] = 8'd14;
        rom[144][21] = -8'd15;
        rom[144][22] = -8'd9;
        rom[144][23] = -8'd5;
        rom[144][24] = 8'd26;
        rom[144][25] = -8'd8;
        rom[144][26] = -8'd36;
        rom[144][27] = 8'd3;
        rom[144][28] = -8'd43;
        rom[144][29] = -8'd4;
        rom[144][30] = -8'd53;
        rom[144][31] = -8'd28;
        rom[145][0] = -8'd25;
        rom[145][1] = -8'd30;
        rom[145][2] = -8'd3;
        rom[145][3] = -8'd6;
        rom[145][4] = -8'd7;
        rom[145][5] = 8'd10;
        rom[145][6] = -8'd13;
        rom[145][7] = -8'd11;
        rom[145][8] = 8'd21;
        rom[145][9] = -8'd26;
        rom[145][10] = 8'd4;
        rom[145][11] = -8'd8;
        rom[145][12] = 8'd5;
        rom[145][13] = -8'd17;
        rom[145][14] = -8'd19;
        rom[145][15] = -8'd17;
        rom[145][16] = -8'd14;
        rom[145][17] = 8'd45;
        rom[145][18] = -8'd58;
        rom[145][19] = 8'd1;
        rom[145][20] = -8'd43;
        rom[145][21] = -8'd66;
        rom[145][22] = 8'd1;
        rom[145][23] = -8'd5;
        rom[145][24] = -8'd13;
        rom[145][25] = 8'd1;
        rom[145][26] = 8'd26;
        rom[145][27] = -8'd34;
        rom[145][28] = -8'd10;
        rom[145][29] = -8'd2;
        rom[145][30] = -8'd2;
        rom[145][31] = 8'd17;
        rom[146][0] = -8'd17;
        rom[146][1] = -8'd27;
        rom[146][2] = 8'd41;
        rom[146][3] = 8'd50;
        rom[146][4] = -8'd13;
        rom[146][5] = 8'd12;
        rom[146][6] = 8'd4;
        rom[146][7] = 8'd2;
        rom[146][8] = 8'd16;
        rom[146][9] = -8'd52;
        rom[146][10] = -8'd24;
        rom[146][11] = 8'd37;
        rom[146][12] = -8'd65;
        rom[146][13] = -8'd56;
        rom[146][14] = -8'd10;
        rom[146][15] = -8'd18;
        rom[146][16] = -8'd39;
        rom[146][17] = -8'd41;
        rom[146][18] = 8'd6;
        rom[146][19] = -8'd37;
        rom[146][20] = -8'd24;
        rom[146][21] = -8'd33;
        rom[146][22] = 8'd44;
        rom[146][23] = -8'd40;
        rom[146][24] = -8'd41;
        rom[146][25] = 8'd20;
        rom[146][26] = -8'd9;
        rom[146][27] = -8'd53;
        rom[146][28] = 8'd30;
        rom[146][29] = 8'd4;
        rom[146][30] = 8'd21;
        rom[146][31] = 8'd29;
        rom[147][0] = 8'd22;
        rom[147][1] = -8'd16;
        rom[147][2] = 8'd8;
        rom[147][3] = 8'd31;
        rom[147][4] = -8'd14;
        rom[147][5] = 8'd11;
        rom[147][6] = 8'd2;
        rom[147][7] = -8'd23;
        rom[147][8] = -8'd26;
        rom[147][9] = 8'd22;
        rom[147][10] = 8'd1;
        rom[147][11] = 8'd10;
        rom[147][12] = -8'd58;
        rom[147][13] = -8'd4;
        rom[147][14] = 8'd4;
        rom[147][15] = 8'd42;
        rom[147][16] = -8'd8;
        rom[147][17] = -8'd4;
        rom[147][18] = 8'd42;
        rom[147][19] = -8'd14;
        rom[147][20] = 8'd28;
        rom[147][21] = 8'd26;
        rom[147][22] = 8'd45;
        rom[147][23] = -8'd55;
        rom[147][24] = -8'd27;
        rom[147][25] = -8'd37;
        rom[147][26] = -8'd5;
        rom[147][27] = 8'd0;
        rom[147][28] = -8'd16;
        rom[147][29] = -8'd12;
        rom[147][30] = 8'd36;
        rom[147][31] = -8'd40;
        rom[148][0] = 8'd40;
        rom[148][1] = 8'd33;
        rom[148][2] = -8'd32;
        rom[148][3] = 8'd13;
        rom[148][4] = 8'd17;
        rom[148][5] = 8'd18;
        rom[148][6] = -8'd5;
        rom[148][7] = -8'd31;
        rom[148][8] = -8'd12;
        rom[148][9] = 8'd12;
        rom[148][10] = 8'd7;
        rom[148][11] = -8'd14;
        rom[148][12] = 8'd5;
        rom[148][13] = -8'd16;
        rom[148][14] = -8'd13;
        rom[148][15] = -8'd27;
        rom[148][16] = -8'd4;
        rom[148][17] = 8'd14;
        rom[148][18] = -8'd15;
        rom[148][19] = -8'd34;
        rom[148][20] = 8'd0;
        rom[148][21] = 8'd20;
        rom[148][22] = -8'd52;
        rom[148][23] = 8'd33;
        rom[148][24] = 8'd28;
        rom[148][25] = 8'd18;
        rom[148][26] = -8'd24;
        rom[148][27] = 8'd15;
        rom[148][28] = -8'd28;
        rom[148][29] = 8'd1;
        rom[148][30] = -8'd57;
        rom[148][31] = -8'd42;
        rom[149][0] = -8'd26;
        rom[149][1] = -8'd22;
        rom[149][2] = -8'd63;
        rom[149][3] = -8'd16;
        rom[149][4] = 8'd6;
        rom[149][5] = -8'd8;
        rom[149][6] = -8'd17;
        rom[149][7] = -8'd1;
        rom[149][8] = 8'd12;
        rom[149][9] = -8'd10;
        rom[149][10] = -8'd9;
        rom[149][11] = -8'd74;
        rom[149][12] = -8'd48;
        rom[149][13] = 8'd21;
        rom[149][14] = 8'd19;
        rom[149][15] = 8'd8;
        rom[149][16] = -8'd5;
        rom[149][17] = -8'd38;
        rom[149][18] = -8'd32;
        rom[149][19] = 8'd6;
        rom[149][20] = -8'd4;
        rom[149][21] = 8'd3;
        rom[149][22] = -8'd18;
        rom[149][23] = 8'd17;
        rom[149][24] = 8'd45;
        rom[149][25] = -8'd15;
        rom[149][26] = -8'd4;
        rom[149][27] = 8'd15;
        rom[149][28] = -8'd15;
        rom[149][29] = -8'd12;
        rom[149][30] = -8'd46;
        rom[149][31] = -8'd24;
        rom[150][0] = -8'd26;
        rom[150][1] = -8'd38;
        rom[150][2] = -8'd5;
        rom[150][3] = 8'd39;
        rom[150][4] = -8'd3;
        rom[150][5] = 8'd21;
        rom[150][6] = -8'd7;
        rom[150][7] = 8'd3;
        rom[150][8] = 8'd12;
        rom[150][9] = 8'd27;
        rom[150][10] = 8'd36;
        rom[150][11] = 8'd19;
        rom[150][12] = -8'd14;
        rom[150][13] = 8'd1;
        rom[150][14] = 8'd1;
        rom[150][15] = 8'd26;
        rom[150][16] = 8'd8;
        rom[150][17] = 8'd27;
        rom[150][18] = 8'd19;
        rom[150][19] = 8'd21;
        rom[150][20] = 8'd10;
        rom[150][21] = -8'd25;
        rom[150][22] = 8'd11;
        rom[150][23] = -8'd2;
        rom[150][24] = -8'd28;
        rom[150][25] = -8'd25;
        rom[150][26] = -8'd21;
        rom[150][27] = -8'd38;
        rom[150][28] = -8'd6;
        rom[150][29] = -8'd3;
        rom[150][30] = -8'd4;
        rom[150][31] = 8'd32;
        rom[151][0] = 8'd2;
        rom[151][1] = 8'd15;
        rom[151][2] = -8'd39;
        rom[151][3] = -8'd19;
        rom[151][4] = 8'd3;
        rom[151][5] = 8'd45;
        rom[151][6] = 8'd2;
        rom[151][7] = -8'd13;
        rom[151][8] = -8'd25;
        rom[151][9] = 8'd4;
        rom[151][10] = -8'd48;
        rom[151][11] = 8'd3;
        rom[151][12] = 8'd20;
        rom[151][13] = -8'd25;
        rom[151][14] = -8'd4;
        rom[151][15] = 8'd19;
        rom[151][16] = 8'd5;
        rom[151][17] = -8'd16;
        rom[151][18] = -8'd22;
        rom[151][19] = -8'd5;
        rom[151][20] = 8'd17;
        rom[151][21] = 8'd1;
        rom[151][22] = -8'd58;
        rom[151][23] = 8'd10;
        rom[151][24] = -8'd35;
        rom[151][25] = -8'd22;
        rom[151][26] = -8'd17;
        rom[151][27] = -8'd2;
        rom[151][28] = 8'd18;
        rom[151][29] = -8'd11;
        rom[151][30] = -8'd12;
        rom[151][31] = 8'd24;
        rom[152][0] = -8'd19;
        rom[152][1] = -8'd27;
        rom[152][2] = -8'd10;
        rom[152][3] = -8'd22;
        rom[152][4] = -8'd92;
        rom[152][5] = 8'd28;
        rom[152][6] = -8'd7;
        rom[152][7] = 8'd7;
        rom[152][8] = 8'd0;
        rom[152][9] = -8'd21;
        rom[152][10] = -8'd5;
        rom[152][11] = -8'd17;
        rom[152][12] = -8'd50;
        rom[152][13] = 8'd43;
        rom[152][14] = 8'd46;
        rom[152][15] = -8'd24;
        rom[152][16] = -8'd2;
        rom[152][17] = -8'd74;
        rom[152][18] = 8'd16;
        rom[152][19] = -8'd35;
        rom[152][20] = 8'd60;
        rom[152][21] = 8'd21;
        rom[152][22] = -8'd34;
        rom[152][23] = -8'd21;
        rom[152][24] = 8'd19;
        rom[152][25] = -8'd21;
        rom[152][26] = -8'd23;
        rom[152][27] = 8'd5;
        rom[152][28] = -8'd13;
        rom[152][29] = -8'd15;
        rom[152][30] = -8'd86;
        rom[152][31] = -8'd13;
        rom[153][0] = -8'd12;
        rom[153][1] = -8'd13;
        rom[153][2] = -8'd24;
        rom[153][3] = -8'd26;
        rom[153][4] = -8'd16;
        rom[153][5] = 8'd63;
        rom[153][6] = 8'd41;
        rom[153][7] = 8'd8;
        rom[153][8] = 8'd22;
        rom[153][9] = 8'd6;
        rom[153][10] = -8'd2;
        rom[153][11] = -8'd25;
        rom[153][12] = -8'd17;
        rom[153][13] = 8'd19;
        rom[153][14] = 8'd11;
        rom[153][15] = 8'd25;
        rom[153][16] = 8'd24;
        rom[153][17] = 8'd26;
        rom[153][18] = -8'd27;
        rom[153][19] = 8'd21;
        rom[153][20] = -8'd17;
        rom[153][21] = 8'd28;
        rom[153][22] = -8'd43;
        rom[153][23] = -8'd46;
        rom[153][24] = 8'd13;
        rom[153][25] = -8'd79;
        rom[153][26] = 8'd12;
        rom[153][27] = -8'd25;
        rom[153][28] = 8'd26;
        rom[153][29] = -8'd2;
        rom[153][30] = -8'd62;
        rom[153][31] = -8'd10;
        rom[154][0] = -8'd48;
        rom[154][1] = -8'd4;
        rom[154][2] = 8'd40;
        rom[154][3] = -8'd34;
        rom[154][4] = 8'd0;
        rom[154][5] = 8'd34;
        rom[154][6] = -8'd23;
        rom[154][7] = -8'd1;
        rom[154][8] = -8'd7;
        rom[154][9] = 8'd14;
        rom[154][10] = -8'd40;
        rom[154][11] = -8'd25;
        rom[154][12] = -8'd24;
        rom[154][13] = -8'd22;
        rom[154][14] = -8'd12;
        rom[154][15] = -8'd19;
        rom[154][16] = 8'd12;
        rom[154][17] = -8'd34;
        rom[154][18] = -8'd46;
        rom[154][19] = 8'd20;
        rom[154][20] = -8'd9;
        rom[154][21] = -8'd8;
        rom[154][22] = -8'd9;
        rom[154][23] = 8'd19;
        rom[154][24] = -8'd10;
        rom[154][25] = -8'd22;
        rom[154][26] = 8'd44;
        rom[154][27] = -8'd35;
        rom[154][28] = 8'd6;
        rom[154][29] = -8'd11;
        rom[154][30] = -8'd8;
        rom[154][31] = -8'd12;
        rom[155][0] = 8'd10;
        rom[155][1] = 8'd0;
        rom[155][2] = -8'd9;
        rom[155][3] = 8'd3;
        rom[155][4] = -8'd1;
        rom[155][5] = -8'd27;
        rom[155][6] = -8'd11;
        rom[155][7] = 8'd1;
        rom[155][8] = -8'd7;
        rom[155][9] = -8'd30;
        rom[155][10] = 8'd0;
        rom[155][11] = 8'd21;
        rom[155][12] = 8'd41;
        rom[155][13] = -8'd8;
        rom[155][14] = -8'd54;
        rom[155][15] = 8'd23;
        rom[155][16] = 8'd6;
        rom[155][17] = -8'd54;
        rom[155][18] = 8'd27;
        rom[155][19] = 8'd4;
        rom[155][20] = -8'd10;
        rom[155][21] = 8'd5;
        rom[155][22] = -8'd45;
        rom[155][23] = -8'd1;
        rom[155][24] = -8'd4;
        rom[155][25] = 8'd25;
        rom[155][26] = -8'd11;
        rom[155][27] = 8'd6;
        rom[155][28] = -8'd5;
        rom[155][29] = 8'd4;
        rom[155][30] = -8'd8;
        rom[155][31] = 8'd37;
        rom[156][0] = -8'd13;
        rom[156][1] = 8'd7;
        rom[156][2] = 8'd23;
        rom[156][3] = 8'd3;
        rom[156][4] = 8'd17;
        rom[156][5] = -8'd24;
        rom[156][6] = 8'd18;
        rom[156][7] = 8'd18;
        rom[156][8] = 8'd19;
        rom[156][9] = 8'd14;
        rom[156][10] = -8'd20;
        rom[156][11] = 8'd0;
        rom[156][12] = 8'd6;
        rom[156][13] = -8'd42;
        rom[156][14] = -8'd15;
        rom[156][15] = -8'd15;
        rom[156][16] = -8'd16;
        rom[156][17] = -8'd12;
        rom[156][18] = -8'd1;
        rom[156][19] = 8'd7;
        rom[156][20] = -8'd47;
        rom[156][21] = 8'd7;
        rom[156][22] = -8'd8;
        rom[156][23] = 8'd6;
        rom[156][24] = 8'd28;
        rom[156][25] = 8'd24;
        rom[156][26] = -8'd9;
        rom[156][27] = -8'd46;
        rom[156][28] = -8'd20;
        rom[156][29] = -8'd17;
        rom[156][30] = 8'd7;
        rom[156][31] = -8'd35;
        rom[157][0] = -8'd22;
        rom[157][1] = -8'd15;
        rom[157][2] = -8'd36;
        rom[157][3] = -8'd4;
        rom[157][4] = 8'd3;
        rom[157][5] = 8'd50;
        rom[157][6] = 8'd57;
        rom[157][7] = -8'd77;
        rom[157][8] = 8'd12;
        rom[157][9] = 8'd38;
        rom[157][10] = 8'd2;
        rom[157][11] = -8'd24;
        rom[157][12] = -8'd34;
        rom[157][13] = 8'd36;
        rom[157][14] = -8'd20;
        rom[157][15] = -8'd15;
        rom[157][16] = 8'd47;
        rom[157][17] = 8'd25;
        rom[157][18] = 8'd11;
        rom[157][19] = 8'd12;
        rom[157][20] = 8'd15;
        rom[157][21] = 8'd13;
        rom[157][22] = -8'd24;
        rom[157][23] = 8'd8;
        rom[157][24] = -8'd37;
        rom[157][25] = -8'd10;
        rom[157][26] = -8'd24;
        rom[157][27] = -8'd10;
        rom[157][28] = 8'd19;
        rom[157][29] = -8'd4;
        rom[157][30] = -8'd10;
        rom[157][31] = -8'd64;
        rom[158][0] = -8'd35;
        rom[158][1] = 8'd52;
        rom[158][2] = -8'd18;
        rom[158][3] = -8'd46;
        rom[158][4] = -8'd10;
        rom[158][5] = 8'd11;
        rom[158][6] = 8'd9;
        rom[158][7] = -8'd8;
        rom[158][8] = 8'd18;
        rom[158][9] = -8'd46;
        rom[158][10] = -8'd13;
        rom[158][11] = 8'd17;
        rom[158][12] = 8'd55;
        rom[158][13] = -8'd21;
        rom[158][14] = 8'd1;
        rom[158][15] = 8'd44;
        rom[158][16] = 8'd22;
        rom[158][17] = 8'd36;
        rom[158][18] = 8'd21;
        rom[158][19] = -8'd6;
        rom[158][20] = -8'd13;
        rom[158][21] = -8'd15;
        rom[158][22] = -8'd34;
        rom[158][23] = -8'd6;
        rom[158][24] = 8'd35;
        rom[158][25] = 8'd49;
        rom[158][26] = 8'd4;
        rom[158][27] = -8'd11;
        rom[158][28] = -8'd18;
        rom[158][29] = -8'd8;
        rom[158][30] = -8'd89;
        rom[158][31] = -8'd43;
        rom[159][0] = -8'd27;
        rom[159][1] = -8'd15;
        rom[159][2] = 8'd28;
        rom[159][3] = 8'd30;
        rom[159][4] = 8'd41;
        rom[159][5] = -8'd41;
        rom[159][6] = -8'd1;
        rom[159][7] = 8'd13;
        rom[159][8] = 8'd21;
        rom[159][9] = -8'd79;
        rom[159][10] = -8'd7;
        rom[159][11] = -8'd9;
        rom[159][12] = 8'd30;
        rom[159][13] = -8'd22;
        rom[159][14] = -8'd37;
        rom[159][15] = 8'd15;
        rom[159][16] = -8'd18;
        rom[159][17] = -8'd7;
        rom[159][18] = 8'd38;
        rom[159][19] = -8'd27;
        rom[159][20] = -8'd14;
        rom[159][21] = -8'd54;
        rom[159][22] = -8'd3;
        rom[159][23] = -8'd25;
        rom[159][24] = 8'd14;
        rom[159][25] = -8'd44;
        rom[159][26] = -8'd34;
        rom[159][27] = -8'd16;
        rom[159][28] = -8'd20;
        rom[159][29] = -8'd13;
        rom[159][30] = 8'd36;
        rom[159][31] = -8'd3;
        rom[160][0] = 8'd28;
        rom[160][1] = -8'd24;
        rom[160][2] = -8'd54;
        rom[160][3] = -8'd56;
        rom[160][4] = 8'd17;
        rom[160][5] = 8'd13;
        rom[160][6] = 8'd22;
        rom[160][7] = -8'd56;
        rom[160][8] = -8'd35;
        rom[160][9] = -8'd7;
        rom[160][10] = 8'd6;
        rom[160][11] = 8'd1;
        rom[160][12] = 8'd0;
        rom[160][13] = 8'd22;
        rom[160][14] = 8'd2;
        rom[160][15] = -8'd9;
        rom[160][16] = -8'd53;
        rom[160][17] = -8'd14;
        rom[160][18] = -8'd6;
        rom[160][19] = -8'd9;
        rom[160][20] = -8'd41;
        rom[160][21] = -8'd9;
        rom[160][22] = 8'd12;
        rom[160][23] = 8'd43;
        rom[160][24] = 8'd1;
        rom[160][25] = -8'd2;
        rom[160][26] = -8'd24;
        rom[160][27] = 8'd5;
        rom[160][28] = 8'd24;
        rom[160][29] = -8'd1;
        rom[160][30] = 8'd14;
        rom[160][31] = 8'd33;
        rom[161][0] = -8'd17;
        rom[161][1] = 8'd41;
        rom[161][2] = 8'd21;
        rom[161][3] = -8'd39;
        rom[161][4] = -8'd52;
        rom[161][5] = -8'd11;
        rom[161][6] = 8'd1;
        rom[161][7] = 8'd41;
        rom[161][8] = 8'd20;
        rom[161][9] = 8'd24;
        rom[161][10] = 8'd6;
        rom[161][11] = 8'd7;
        rom[161][12] = 8'd48;
        rom[161][13] = -8'd34;
        rom[161][14] = 8'd13;
        rom[161][15] = -8'd14;
        rom[161][16] = 8'd43;
        rom[161][17] = -8'd20;
        rom[161][18] = 8'd39;
        rom[161][19] = -8'd2;
        rom[161][20] = 8'd3;
        rom[161][21] = -8'd4;
        rom[161][22] = -8'd1;
        rom[161][23] = -8'd45;
        rom[161][24] = 8'd53;
        rom[161][25] = 8'd36;
        rom[161][26] = -8'd22;
        rom[161][27] = 8'd7;
        rom[161][28] = -8'd2;
        rom[161][29] = -8'd1;
        rom[161][30] = -8'd66;
        rom[161][31] = 8'd15;
        rom[162][0] = 8'd3;
        rom[162][1] = -8'd62;
        rom[162][2] = -8'd101;
        rom[162][3] = 8'd9;
        rom[162][4] = 8'd4;
        rom[162][5] = 8'd19;
        rom[162][6] = 8'd10;
        rom[162][7] = -8'd56;
        rom[162][8] = -8'd35;
        rom[162][9] = -8'd10;
        rom[162][10] = 8'd2;
        rom[162][11] = -8'd37;
        rom[162][12] = 8'd19;
        rom[162][13] = -8'd12;
        rom[162][14] = -8'd58;
        rom[162][15] = -8'd40;
        rom[162][16] = -8'd11;
        rom[162][17] = 8'd11;
        rom[162][18] = -8'd37;
        rom[162][19] = -8'd44;
        rom[162][20] = -8'd21;
        rom[162][21] = 8'd28;
        rom[162][22] = 8'd1;
        rom[162][23] = 8'd30;
        rom[162][24] = 8'd1;
        rom[162][25] = -8'd91;
        rom[162][26] = 8'd1;
        rom[162][27] = -8'd7;
        rom[162][28] = -8'd13;
        rom[162][29] = 8'd10;
        rom[162][30] = 8'd4;
        rom[162][31] = 8'd15;
        rom[163][0] = 8'd6;
        rom[163][1] = -8'd26;
        rom[163][2] = -8'd21;
        rom[163][3] = 8'd19;
        rom[163][4] = -8'd9;
        rom[163][5] = 8'd16;
        rom[163][6] = 8'd27;
        rom[163][7] = -8'd12;
        rom[163][8] = 8'd4;
        rom[163][9] = -8'd41;
        rom[163][10] = -8'd47;
        rom[163][11] = -8'd14;
        rom[163][12] = -8'd21;
        rom[163][13] = -8'd11;
        rom[163][14] = -8'd26;
        rom[163][15] = 8'd16;
        rom[163][16] = 8'd7;
        rom[163][17] = 8'd9;
        rom[163][18] = 8'd0;
        rom[163][19] = -8'd12;
        rom[163][20] = 8'd28;
        rom[163][21] = -8'd39;
        rom[163][22] = -8'd12;
        rom[163][23] = -8'd6;
        rom[163][24] = 8'd17;
        rom[163][25] = 8'd26;
        rom[163][26] = -8'd3;
        rom[163][27] = 8'd7;
        rom[163][28] = -8'd32;
        rom[163][29] = -8'd7;
        rom[163][30] = 8'd3;
        rom[163][31] = -8'd19;
        rom[164][0] = -8'd59;
        rom[164][1] = 8'd13;
        rom[164][2] = 8'd22;
        rom[164][3] = 8'd20;
        rom[164][4] = -8'd33;
        rom[164][5] = -8'd4;
        rom[164][6] = 8'd18;
        rom[164][7] = 8'd50;
        rom[164][8] = 8'd8;
        rom[164][9] = 8'd1;
        rom[164][10] = 8'd0;
        rom[164][11] = -8'd4;
        rom[164][12] = -8'd16;
        rom[164][13] = -8'd19;
        rom[164][14] = 8'd51;
        rom[164][15] = 8'd33;
        rom[164][16] = 8'd17;
        rom[164][17] = -8'd8;
        rom[164][18] = 8'd8;
        rom[164][19] = -8'd13;
        rom[164][20] = 8'd24;
        rom[164][21] = 8'd14;
        rom[164][22] = -8'd88;
        rom[164][23] = 8'd16;
        rom[164][24] = 8'd34;
        rom[164][25] = -8'd23;
        rom[164][26] = -8'd23;
        rom[164][27] = -8'd30;
        rom[164][28] = -8'd40;
        rom[164][29] = 8'd8;
        rom[164][30] = -8'd8;
        rom[164][31] = 8'd30;
        rom[165][0] = 8'd43;
        rom[165][1] = -8'd17;
        rom[165][2] = -8'd50;
        rom[165][3] = -8'd37;
        rom[165][4] = -8'd4;
        rom[165][5] = 8'd19;
        rom[165][6] = 8'd18;
        rom[165][7] = -8'd56;
        rom[165][8] = 8'd25;
        rom[165][9] = 8'd3;
        rom[165][10] = -8'd17;
        rom[165][11] = 8'd13;
        rom[165][12] = -8'd4;
        rom[165][13] = 8'd53;
        rom[165][14] = 8'd13;
        rom[165][15] = -8'd23;
        rom[165][16] = 8'd30;
        rom[165][17] = 8'd28;
        rom[165][18] = -8'd40;
        rom[165][19] = 8'd3;
        rom[165][20] = -8'd30;
        rom[165][21] = 8'd33;
        rom[165][22] = -8'd6;
        rom[165][23] = 8'd20;
        rom[165][24] = -8'd18;
        rom[165][25] = -8'd56;
        rom[165][26] = -8'd17;
        rom[165][27] = 8'd22;
        rom[165][28] = -8'd7;
        rom[165][29] = -8'd9;
        rom[165][30] = 8'd0;
        rom[165][31] = 8'd0;
        rom[166][0] = -8'd3;
        rom[166][1] = 8'd21;
        rom[166][2] = 8'd22;
        rom[166][3] = -8'd20;
        rom[166][4] = -8'd2;
        rom[166][5] = -8'd1;
        rom[166][6] = -8'd10;
        rom[166][7] = -8'd18;
        rom[166][8] = -8'd14;
        rom[166][9] = -8'd25;
        rom[166][10] = -8'd47;
        rom[166][11] = -8'd10;
        rom[166][12] = 8'd20;
        rom[166][13] = 8'd9;
        rom[166][14] = 8'd1;
        rom[166][15] = -8'd24;
        rom[166][16] = 8'd10;
        rom[166][17] = 8'd8;
        rom[166][18] = -8'd41;
        rom[166][19] = 8'd13;
        rom[166][20] = -8'd10;
        rom[166][21] = 8'd2;
        rom[166][22] = 8'd8;
        rom[166][23] = -8'd36;
        rom[166][24] = 8'd3;
        rom[166][25] = -8'd55;
        rom[166][26] = -8'd3;
        rom[166][27] = -8'd36;
        rom[166][28] = 8'd36;
        rom[166][29] = -8'd2;
        rom[166][30] = -8'd19;
        rom[166][31] = 8'd24;
        rom[167][0] = -8'd15;
        rom[167][1] = 8'd12;
        rom[167][2] = 8'd34;
        rom[167][3] = -8'd3;
        rom[167][4] = 8'd22;
        rom[167][5] = -8'd54;
        rom[167][6] = -8'd26;
        rom[167][7] = -8'd3;
        rom[167][8] = 8'd32;
        rom[167][9] = 8'd0;
        rom[167][10] = -8'd2;
        rom[167][11] = -8'd7;
        rom[167][12] = 8'd27;
        rom[167][13] = 8'd4;
        rom[167][14] = -8'd45;
        rom[167][15] = 8'd22;
        rom[167][16] = -8'd6;
        rom[167][17] = -8'd9;
        rom[167][18] = 8'd11;
        rom[167][19] = -8'd11;
        rom[167][20] = -8'd21;
        rom[167][21] = -8'd12;
        rom[167][22] = -8'd10;
        rom[167][23] = -8'd22;
        rom[167][24] = 8'd16;
        rom[167][25] = 8'd21;
        rom[167][26] = 8'd41;
        rom[167][27] = 8'd4;
        rom[167][28] = 8'd11;
        rom[167][29] = -8'd5;
        rom[167][30] = -8'd8;
        rom[167][31] = 8'd10;
        rom[168][0] = -8'd10;
        rom[168][1] = -8'd30;
        rom[168][2] = -8'd7;
        rom[168][3] = 8'd13;
        rom[168][4] = -8'd11;
        rom[168][5] = -8'd32;
        rom[168][6] = 8'd36;
        rom[168][7] = -8'd25;
        rom[168][8] = 8'd13;
        rom[168][9] = -8'd8;
        rom[168][10] = 8'd18;
        rom[168][11] = 8'd9;
        rom[168][12] = 8'd8;
        rom[168][13] = -8'd33;
        rom[168][14] = 8'd31;
        rom[168][15] = -8'd11;
        rom[168][16] = -8'd49;
        rom[168][17] = 8'd21;
        rom[168][18] = 8'd1;
        rom[168][19] = -8'd35;
        rom[168][20] = -8'd36;
        rom[168][21] = -8'd21;
        rom[168][22] = 8'd5;
        rom[168][23] = 8'd14;
        rom[168][24] = 8'd33;
        rom[168][25] = -8'd8;
        rom[168][26] = -8'd11;
        rom[168][27] = -8'd15;
        rom[168][28] = -8'd50;
        rom[168][29] = -8'd8;
        rom[168][30] = -8'd39;
        rom[168][31] = 8'd1;
        rom[169][0] = -8'd7;
        rom[169][1] = -8'd23;
        rom[169][2] = 8'd11;
        rom[169][3] = -8'd1;
        rom[169][4] = 8'd9;
        rom[169][5] = -8'd3;
        rom[169][6] = 8'd18;
        rom[169][7] = 8'd16;
        rom[169][8] = -8'd57;
        rom[169][9] = 8'd30;
        rom[169][10] = 8'd2;
        rom[169][11] = -8'd30;
        rom[169][12] = 8'd4;
        rom[169][13] = -8'd25;
        rom[169][14] = -8'd31;
        rom[169][15] = 8'd36;
        rom[169][16] = 8'd1;
        rom[169][17] = -8'd58;
        rom[169][18] = -8'd21;
        rom[169][19] = -8'd19;
        rom[169][20] = 8'd24;
        rom[169][21] = -8'd14;
        rom[169][22] = 8'd1;
        rom[169][23] = 8'd18;
        rom[169][24] = 8'd18;
        rom[169][25] = -8'd27;
        rom[169][26] = 8'd20;
        rom[169][27] = 8'd3;
        rom[169][28] = 8'd3;
        rom[169][29] = -8'd5;
        rom[169][30] = -8'd1;
        rom[169][31] = 8'd44;
        rom[170][0] = 8'd6;
        rom[170][1] = -8'd26;
        rom[170][2] = -8'd36;
        rom[170][3] = -8'd17;
        rom[170][4] = 8'd15;
        rom[170][5] = 8'd25;
        rom[170][6] = 8'd3;
        rom[170][7] = -8'd15;
        rom[170][8] = -8'd11;
        rom[170][9] = 8'd22;
        rom[170][10] = 8'd1;
        rom[170][11] = -8'd3;
        rom[170][12] = -8'd21;
        rom[170][13] = -8'd31;
        rom[170][14] = -8'd10;
        rom[170][15] = 8'd16;
        rom[170][16] = 8'd2;
        rom[170][17] = 8'd52;
        rom[170][18] = -8'd46;
        rom[170][19] = -8'd13;
        rom[170][20] = -8'd19;
        rom[170][21] = 8'd18;
        rom[170][22] = 8'd16;
        rom[170][23] = -8'd30;
        rom[170][24] = 8'd13;
        rom[170][25] = -8'd11;
        rom[170][26] = -8'd4;
        rom[170][27] = -8'd32;
        rom[170][28] = -8'd1;
        rom[170][29] = -8'd15;
        rom[170][30] = 8'd48;
        rom[170][31] = -8'd27;
        rom[171][0] = 8'd33;
        rom[171][1] = 8'd3;
        rom[171][2] = -8'd11;
        rom[171][3] = -8'd26;
        rom[171][4] = -8'd27;
        rom[171][5] = 8'd5;
        rom[171][6] = -8'd14;
        rom[171][7] = -8'd57;
        rom[171][8] = 8'd19;
        rom[171][9] = 8'd10;
        rom[171][10] = -8'd16;
        rom[171][11] = -8'd27;
        rom[171][12] = -8'd61;
        rom[171][13] = 8'd19;
        rom[171][14] = 8'd0;
        rom[171][15] = 8'd5;
        rom[171][16] = 8'd39;
        rom[171][17] = -8'd8;
        rom[171][18] = 8'd22;
        rom[171][19] = -8'd1;
        rom[171][20] = 8'd31;
        rom[171][21] = 8'd37;
        rom[171][22] = -8'd19;
        rom[171][23] = -8'd42;
        rom[171][24] = 8'd16;
        rom[171][25] = -8'd1;
        rom[171][26] = 8'd16;
        rom[171][27] = 8'd16;
        rom[171][28] = 8'd11;
        rom[171][29] = -8'd14;
        rom[171][30] = -8'd16;
        rom[171][31] = -8'd48;
        rom[172][0] = 8'd59;
        rom[172][1] = -8'd1;
        rom[172][2] = -8'd24;
        rom[172][3] = -8'd13;
        rom[172][4] = -8'd17;
        rom[172][5] = -8'd19;
        rom[172][6] = 8'd3;
        rom[172][7] = -8'd35;
        rom[172][8] = -8'd3;
        rom[172][9] = -8'd4;
        rom[172][10] = 8'd45;
        rom[172][11] = 8'd39;
        rom[172][12] = 8'd12;
        rom[172][13] = -8'd2;
        rom[172][14] = -8'd23;
        rom[172][15] = 8'd33;
        rom[172][16] = 8'd19;
        rom[172][17] = -8'd1;
        rom[172][18] = 8'd8;
        rom[172][19] = 8'd12;
        rom[172][20] = -8'd16;
        rom[172][21] = 8'd14;
        rom[172][22] = 8'd12;
        rom[172][23] = 8'd44;
        rom[172][24] = 8'd13;
        rom[172][25] = 8'd19;
        rom[172][26] = -8'd9;
        rom[172][27] = 8'd13;
        rom[172][28] = -8'd45;
        rom[172][29] = -8'd17;
        rom[172][30] = -8'd27;
        rom[172][31] = 8'd16;
        rom[173][0] = 8'd23;
        rom[173][1] = -8'd41;
        rom[173][2] = 8'd0;
        rom[173][3] = -8'd17;
        rom[173][4] = 8'd2;
        rom[173][5] = 8'd4;
        rom[173][6] = -8'd28;
        rom[173][7] = -8'd14;
        rom[173][8] = -8'd18;
        rom[173][9] = -8'd7;
        rom[173][10] = 8'd0;
        rom[173][11] = 8'd31;
        rom[173][12] = -8'd53;
        rom[173][13] = -8'd29;
        rom[173][14] = -8'd27;
        rom[173][15] = 8'd18;
        rom[173][16] = -8'd11;
        rom[173][17] = -8'd35;
        rom[173][18] = -8'd11;
        rom[173][19] = 8'd28;
        rom[173][20] = -8'd15;
        rom[173][21] = -8'd1;
        rom[173][22] = -8'd5;
        rom[173][23] = 8'd12;
        rom[173][24] = -8'd12;
        rom[173][25] = 8'd3;
        rom[173][26] = 8'd6;
        rom[173][27] = 8'd51;
        rom[173][28] = -8'd52;
        rom[173][29] = 8'd11;
        rom[173][30] = 8'd22;
        rom[173][31] = -8'd30;
        rom[174][0] = -8'd18;
        rom[174][1] = -8'd5;
        rom[174][2] = 8'd30;
        rom[174][3] = -8'd3;
        rom[174][4] = 8'd14;
        rom[174][5] = -8'd2;
        rom[174][6] = -8'd11;
        rom[174][7] = 8'd11;
        rom[174][8] = 8'd9;
        rom[174][9] = 8'd5;
        rom[174][10] = 8'd25;
        rom[174][11] = -8'd30;
        rom[174][12] = 8'd4;
        rom[174][13] = -8'd1;
        rom[174][14] = -8'd13;
        rom[174][15] = 8'd18;
        rom[174][16] = -8'd16;
        rom[174][17] = -8'd61;
        rom[174][18] = 8'd32;
        rom[174][19] = -8'd1;
        rom[174][20] = -8'd16;
        rom[174][21] = -8'd27;
        rom[174][22] = -8'd13;
        rom[174][23] = -8'd7;
        rom[174][24] = 8'd2;
        rom[174][25] = 8'd20;
        rom[174][26] = 8'd4;
        rom[174][27] = -8'd6;
        rom[174][28] = 8'd11;
        rom[174][29] = -8'd7;
        rom[174][30] = 8'd1;
        rom[174][31] = 8'd12;
        rom[175][0] = 8'd16;
        rom[175][1] = -8'd6;
        rom[175][2] = 8'd9;
        rom[175][3] = 8'd4;
        rom[175][4] = -8'd16;
        rom[175][5] = -8'd38;
        rom[175][6] = 8'd18;
        rom[175][7] = 8'd31;
        rom[175][8] = -8'd42;
        rom[175][9] = -8'd55;
        rom[175][10] = -8'd46;
        rom[175][11] = 8'd6;
        rom[175][12] = 8'd8;
        rom[175][13] = -8'd3;
        rom[175][14] = 8'd5;
        rom[175][15] = 8'd8;
        rom[175][16] = -8'd29;
        rom[175][17] = 8'd9;
        rom[175][18] = 8'd2;
        rom[175][19] = 8'd12;
        rom[175][20] = -8'd14;
        rom[175][21] = -8'd14;
        rom[175][22] = 8'd18;
        rom[175][23] = -8'd26;
        rom[175][24] = 8'd15;
        rom[175][25] = -8'd18;
        rom[175][26] = -8'd42;
        rom[175][27] = 8'd0;
        rom[175][28] = -8'd39;
        rom[175][29] = 8'd4;
        rom[175][30] = 8'd3;
        rom[175][31] = 8'd33;
        rom[176][0] = 8'd5;
        rom[176][1] = -8'd10;
        rom[176][2] = 8'd18;
        rom[176][3] = 8'd1;
        rom[176][4] = -8'd21;
        rom[176][5] = 8'd10;
        rom[176][6] = -8'd20;
        rom[176][7] = -8'd37;
        rom[176][8] = 8'd15;
        rom[176][9] = -8'd15;
        rom[176][10] = 8'd3;
        rom[176][11] = -8'd14;
        rom[176][12] = 8'd6;
        rom[176][13] = -8'd29;
        rom[176][14] = -8'd22;
        rom[176][15] = -8'd17;
        rom[176][16] = 8'd32;
        rom[176][17] = 8'd21;
        rom[176][18] = 8'd16;
        rom[176][19] = -8'd64;
        rom[176][20] = -8'd22;
        rom[176][21] = -8'd12;
        rom[176][22] = 8'd7;
        rom[176][23] = 8'd58;
        rom[176][24] = 8'd33;
        rom[176][25] = -8'd17;
        rom[176][26] = -8'd3;
        rom[176][27] = -8'd16;
        rom[176][28] = -8'd32;
        rom[176][29] = 8'd3;
        rom[176][30] = -8'd11;
        rom[176][31] = -8'd6;
        rom[177][0] = 8'd47;
        rom[177][1] = -8'd44;
        rom[177][2] = -8'd18;
        rom[177][3] = 8'd31;
        rom[177][4] = -8'd15;
        rom[177][5] = 8'd23;
        rom[177][6] = -8'd20;
        rom[177][7] = -8'd10;
        rom[177][8] = 8'd16;
        rom[177][9] = -8'd11;
        rom[177][10] = -8'd2;
        rom[177][11] = 8'd8;
        rom[177][12] = 8'd8;
        rom[177][13] = 8'd50;
        rom[177][14] = -8'd20;
        rom[177][15] = 8'd7;
        rom[177][16] = -8'd62;
        rom[177][17] = 8'd9;
        rom[177][18] = -8'd24;
        rom[177][19] = 8'd15;
        rom[177][20] = 8'd1;
        rom[177][21] = -8'd12;
        rom[177][22] = 8'd0;
        rom[177][23] = -8'd3;
        rom[177][24] = -8'd3;
        rom[177][25] = -8'd39;
        rom[177][26] = 8'd25;
        rom[177][27] = 8'd12;
        rom[177][28] = 8'd4;
        rom[177][29] = -8'd17;
        rom[177][30] = -8'd17;
        rom[177][31] = 8'd8;
        rom[178][0] = -8'd3;
        rom[178][1] = -8'd26;
        rom[178][2] = 8'd8;
        rom[178][3] = 8'd40;
        rom[178][4] = -8'd12;
        rom[178][5] = -8'd9;
        rom[178][6] = 8'd29;
        rom[178][7] = 8'd28;
        rom[178][8] = -8'd40;
        rom[178][9] = -8'd35;
        rom[178][10] = -8'd35;
        rom[178][11] = 8'd22;
        rom[178][12] = -8'd21;
        rom[178][13] = -8'd29;
        rom[178][14] = 8'd10;
        rom[178][15] = -8'd26;
        rom[178][16] = -8'd123;
        rom[178][17] = 8'd21;
        rom[178][18] = -8'd19;
        rom[178][19] = -8'd5;
        rom[178][20] = 8'd3;
        rom[178][21] = -8'd19;
        rom[178][22] = 8'd32;
        rom[178][23] = 8'd13;
        rom[178][24] = -8'd18;
        rom[178][25] = 8'd13;
        rom[178][26] = -8'd16;
        rom[178][27] = -8'd48;
        rom[178][28] = -8'd11;
        rom[178][29] = -8'd5;
        rom[178][30] = 8'd29;
        rom[178][31] = 8'd12;
        rom[179][0] = -8'd20;
        rom[179][1] = 8'd20;
        rom[179][2] = 8'd35;
        rom[179][3] = 8'd1;
        rom[179][4] = 8'd26;
        rom[179][5] = 8'd22;
        rom[179][6] = -8'd6;
        rom[179][7] = -8'd62;
        rom[179][8] = -8'd19;
        rom[179][9] = 8'd24;
        rom[179][10] = 8'd35;
        rom[179][11] = 8'd19;
        rom[179][12] = -8'd44;
        rom[179][13] = -8'd28;
        rom[179][14] = -8'd2;
        rom[179][15] = 8'd31;
        rom[179][16] = -8'd3;
        rom[179][17] = 8'd12;
        rom[179][18] = 8'd42;
        rom[179][19] = 8'd1;
        rom[179][20] = 8'd27;
        rom[179][21] = -8'd7;
        rom[179][22] = 8'd17;
        rom[179][23] = 8'd27;
        rom[179][24] = -8'd4;
        rom[179][25] = -8'd8;
        rom[179][26] = -8'd18;
        rom[179][27] = -8'd8;
        rom[179][28] = 8'd13;
        rom[179][29] = -8'd4;
        rom[179][30] = 8'd3;
        rom[179][31] = -8'd43;
        rom[180][0] = 8'd30;
        rom[180][1] = 8'd44;
        rom[180][2] = -8'd26;
        rom[180][3] = 8'd14;
        rom[180][4] = 8'd27;
        rom[180][5] = 8'd28;
        rom[180][6] = 8'd29;
        rom[180][7] = -8'd80;
        rom[180][8] = 8'd40;
        rom[180][9] = 8'd8;
        rom[180][10] = 8'd42;
        rom[180][11] = -8'd30;
        rom[180][12] = 8'd6;
        rom[180][13] = 8'd14;
        rom[180][14] = -8'd10;
        rom[180][15] = 8'd15;
        rom[180][16] = -8'd7;
        rom[180][17] = -8'd3;
        rom[180][18] = -8'd7;
        rom[180][19] = -8'd31;
        rom[180][20] = 8'd11;
        rom[180][21] = 8'd10;
        rom[180][22] = -8'd39;
        rom[180][23] = -8'd4;
        rom[180][24] = 8'd15;
        rom[180][25] = 8'd38;
        rom[180][26] = -8'd19;
        rom[180][27] = 8'd8;
        rom[180][28] = -8'd19;
        rom[180][29] = 8'd2;
        rom[180][30] = -8'd58;
        rom[180][31] = -8'd30;
        rom[181][0] = -8'd10;
        rom[181][1] = -8'd40;
        rom[181][2] = 8'd3;
        rom[181][3] = -8'd14;
        rom[181][4] = 8'd29;
        rom[181][5] = -8'd11;
        rom[181][6] = 8'd30;
        rom[181][7] = -8'd32;
        rom[181][8] = 8'd23;
        rom[181][9] = -8'd4;
        rom[181][10] = -8'd24;
        rom[181][11] = -8'd23;
        rom[181][12] = -8'd6;
        rom[181][13] = -8'd16;
        rom[181][14] = 8'd30;
        rom[181][15] = 8'd20;
        rom[181][16] = 8'd4;
        rom[181][17] = -8'd48;
        rom[181][18] = -8'd35;
        rom[181][19] = -8'd11;
        rom[181][20] = -8'd3;
        rom[181][21] = -8'd2;
        rom[181][22] = -8'd13;
        rom[181][23] = -8'd6;
        rom[181][24] = 8'd17;
        rom[181][25] = -8'd37;
        rom[181][26] = -8'd12;
        rom[181][27] = 8'd32;
        rom[181][28] = -8'd32;
        rom[181][29] = -8'd7;
        rom[181][30] = -8'd23;
        rom[181][31] = -8'd9;
        rom[182][0] = -8'd66;
        rom[182][1] = -8'd47;
        rom[182][2] = 8'd29;
        rom[182][3] = 8'd26;
        rom[182][4] = -8'd16;
        rom[182][5] = 8'd2;
        rom[182][6] = -8'd19;
        rom[182][7] = 8'd34;
        rom[182][8] = 8'd23;
        rom[182][9] = 8'd7;
        rom[182][10] = 8'd38;
        rom[182][11] = 8'd21;
        rom[182][12] = -8'd32;
        rom[182][13] = 8'd19;
        rom[182][14] = -8'd14;
        rom[182][15] = 8'd6;
        rom[182][16] = 8'd1;
        rom[182][17] = -8'd25;
        rom[182][18] = 8'd20;
        rom[182][19] = 8'd26;
        rom[182][20] = 8'd4;
        rom[182][21] = -8'd4;
        rom[182][22] = 8'd9;
        rom[182][23] = -8'd8;
        rom[182][24] = -8'd23;
        rom[182][25] = -8'd48;
        rom[182][26] = 8'd26;
        rom[182][27] = -8'd8;
        rom[182][28] = 8'd29;
        rom[182][29] = 8'd4;
        rom[182][30] = 8'd11;
        rom[182][31] = -8'd7;
        rom[183][0] = 8'd33;
        rom[183][1] = 8'd51;
        rom[183][2] = -8'd10;
        rom[183][3] = 8'd13;
        rom[183][4] = -8'd10;
        rom[183][5] = -8'd22;
        rom[183][6] = -8'd9;
        rom[183][7] = 8'd5;
        rom[183][8] = 8'd7;
        rom[183][9] = -8'd3;
        rom[183][10] = -8'd7;
        rom[183][11] = -8'd14;
        rom[183][12] = 8'd21;
        rom[183][13] = 8'd0;
        rom[183][14] = -8'd16;
        rom[183][15] = 8'd8;
        rom[183][16] = -8'd32;
        rom[183][17] = -8'd18;
        rom[183][18] = -8'd17;
        rom[183][19] = 8'd7;
        rom[183][20] = -8'd11;
        rom[183][21] = 8'd13;
        rom[183][22] = -8'd59;
        rom[183][23] = -8'd50;
        rom[183][24] = -8'd12;
        rom[183][25] = 8'd20;
        rom[183][26] = 8'd0;
        rom[183][27] = 8'd2;
        rom[183][28] = 8'd29;
        rom[183][29] = -8'd11;
        rom[183][30] = -8'd15;
        rom[183][31] = 8'd7;
        rom[184][0] = 8'd5;
        rom[184][1] = -8'd5;
        rom[184][2] = 8'd12;
        rom[184][3] = -8'd60;
        rom[184][4] = -8'd83;
        rom[184][5] = -8'd19;
        rom[184][6] = -8'd14;
        rom[184][7] = -8'd10;
        rom[184][8] = -8'd12;
        rom[184][9] = -8'd10;
        rom[184][10] = 8'd13;
        rom[184][11] = -8'd8;
        rom[184][12] = -8'd52;
        rom[184][13] = 8'd40;
        rom[184][14] = 8'd48;
        rom[184][15] = -8'd32;
        rom[184][16] = 8'd17;
        rom[184][17] = -8'd18;
        rom[184][18] = -8'd9;
        rom[184][19] = -8'd13;
        rom[184][20] = 8'd24;
        rom[184][21] = -8'd18;
        rom[184][22] = -8'd44;
        rom[184][23] = -8'd5;
        rom[184][24] = 8'd15;
        rom[184][25] = 8'd55;
        rom[184][26] = -8'd28;
        rom[184][27] = 8'd8;
        rom[184][28] = -8'd61;
        rom[184][29] = -8'd10;
        rom[184][30] = -8'd55;
        rom[184][31] = -8'd36;
        rom[185][0] = -8'd33;
        rom[185][1] = -8'd5;
        rom[185][2] = 8'd27;
        rom[185][3] = -8'd26;
        rom[185][4] = -8'd22;
        rom[185][5] = 8'd38;
        rom[185][6] = 8'd44;
        rom[185][7] = 8'd21;
        rom[185][8] = 8'd27;
        rom[185][9] = 8'd11;
        rom[185][10] = -8'd5;
        rom[185][11] = -8'd9;
        rom[185][12] = 8'd1;
        rom[185][13] = 8'd2;
        rom[185][14] = 8'd15;
        rom[185][15] = 8'd17;
        rom[185][16] = 8'd31;
        rom[185][17] = 8'd0;
        rom[185][18] = 8'd26;
        rom[185][19] = 8'd7;
        rom[185][20] = -8'd52;
        rom[185][21] = -8'd14;
        rom[185][22] = -8'd88;
        rom[185][23] = -8'd59;
        rom[185][24] = 8'd16;
        rom[185][25] = -8'd55;
        rom[185][26] = 8'd21;
        rom[185][27] = -8'd11;
        rom[185][28] = -8'd2;
        rom[185][29] = -8'd8;
        rom[185][30] = -8'd25;
        rom[185][31] = -8'd6;
        rom[186][0] = 8'd25;
        rom[186][1] = -8'd13;
        rom[186][2] = -8'd14;
        rom[186][3] = -8'd19;
        rom[186][4] = 8'd26;
        rom[186][5] = 8'd25;
        rom[186][6] = -8'd4;
        rom[186][7] = 8'd11;
        rom[186][8] = -8'd17;
        rom[186][9] = 8'd9;
        rom[186][10] = -8'd27;
        rom[186][11] = 8'd8;
        rom[186][12] = -8'd43;
        rom[186][13] = -8'd15;
        rom[186][14] = 8'd1;
        rom[186][15] = -8'd39;
        rom[186][16] = -8'd19;
        rom[186][17] = -8'd32;
        rom[186][18] = -8'd20;
        rom[186][19] = 8'd18;
        rom[186][20] = -8'd7;
        rom[186][21] = 8'd14;
        rom[186][22] = -8'd13;
        rom[186][23] = 8'd6;
        rom[186][24] = 8'd6;
        rom[186][25] = -8'd19;
        rom[186][26] = 8'd19;
        rom[186][27] = -8'd29;
        rom[186][28] = -8'd5;
        rom[186][29] = 8'd7;
        rom[186][30] = -8'd9;
        rom[186][31] = 8'd28;
        rom[187][0] = 8'd13;
        rom[187][1] = -8'd6;
        rom[187][2] = 8'd23;
        rom[187][3] = -8'd7;
        rom[187][4] = 8'd12;
        rom[187][5] = -8'd31;
        rom[187][6] = -8'd8;
        rom[187][7] = -8'd22;
        rom[187][8] = 8'd6;
        rom[187][9] = -8'd2;
        rom[187][10] = 8'd20;
        rom[187][11] = 8'd22;
        rom[187][12] = 8'd8;
        rom[187][13] = -8'd5;
        rom[187][14] = 8'd2;
        rom[187][15] = 8'd39;
        rom[187][16] = 8'd11;
        rom[187][17] = -8'd24;
        rom[187][18] = 8'd21;
        rom[187][19] = 8'd7;
        rom[187][20] = 8'd12;
        rom[187][21] = -8'd26;
        rom[187][22] = -8'd30;
        rom[187][23] = 8'd1;
        rom[187][24] = -8'd2;
        rom[187][25] = 8'd16;
        rom[187][26] = 8'd11;
        rom[187][27] = 8'd3;
        rom[187][28] = 8'd30;
        rom[187][29] = -8'd10;
        rom[187][30] = -8'd5;
        rom[187][31] = 8'd10;
        rom[188][0] = 8'd5;
        rom[188][1] = -8'd1;
        rom[188][2] = -8'd53;
        rom[188][3] = 8'd8;
        rom[188][4] = 8'd11;
        rom[188][5] = 8'd18;
        rom[188][6] = 8'd24;
        rom[188][7] = -8'd16;
        rom[188][8] = -8'd15;
        rom[188][9] = 8'd10;
        rom[188][10] = -8'd5;
        rom[188][11] = 8'd2;
        rom[188][12] = 8'd0;
        rom[188][13] = -8'd5;
        rom[188][14] = -8'd6;
        rom[188][15] = 8'd10;
        rom[188][16] = -8'd24;
        rom[188][17] = -8'd2;
        rom[188][18] = -8'd7;
        rom[188][19] = 8'd3;
        rom[188][20] = 8'd8;
        rom[188][21] = -8'd1;
        rom[188][22] = 8'd4;
        rom[188][23] = 8'd37;
        rom[188][24] = -8'd9;
        rom[188][25] = 8'd33;
        rom[188][26] = 8'd1;
        rom[188][27] = 8'd18;
        rom[188][28] = 8'd0;
        rom[188][29] = -8'd5;
        rom[188][30] = 8'd14;
        rom[188][31] = -8'd26;
        rom[189][0] = -8'd58;
        rom[189][1] = -8'd17;
        rom[189][2] = 8'd15;
        rom[189][3] = -8'd12;
        rom[189][4] = 8'd17;
        rom[189][5] = 8'd23;
        rom[189][6] = 8'd56;
        rom[189][7] = -8'd46;
        rom[189][8] = 8'd31;
        rom[189][9] = 8'd36;
        rom[189][10] = 8'd14;
        rom[189][11] = -8'd8;
        rom[189][12] = -8'd2;
        rom[189][13] = 8'd37;
        rom[189][14] = -8'd8;
        rom[189][15] = 8'd7;
        rom[189][16] = 8'd25;
        rom[189][17] = 8'd3;
        rom[189][18] = -8'd24;
        rom[189][19] = 8'd16;
        rom[189][20] = 8'd17;
        rom[189][21] = 8'd10;
        rom[189][22] = -8'd20;
        rom[189][23] = -8'd22;
        rom[189][24] = -8'd22;
        rom[189][25] = 8'd6;
        rom[189][26] = -8'd12;
        rom[189][27] = -8'd13;
        rom[189][28] = 8'd23;
        rom[189][29] = -8'd1;
        rom[189][30] = 8'd12;
        rom[189][31] = -8'd22;
        rom[190][0] = -8'd53;
        rom[190][1] = 8'd12;
        rom[190][2] = -8'd32;
        rom[190][3] = -8'd45;
        rom[190][4] = 8'd8;
        rom[190][5] = 8'd22;
        rom[190][6] = -8'd13;
        rom[190][7] = -8'd46;
        rom[190][8] = 8'd48;
        rom[190][9] = -8'd1;
        rom[190][10] = -8'd19;
        rom[190][11] = -8'd31;
        rom[190][12] = 8'd18;
        rom[190][13] = -8'd11;
        rom[190][14] = -8'd37;
        rom[190][15] = 8'd33;
        rom[190][16] = 8'd44;
        rom[190][17] = 8'd4;
        rom[190][18] = -8'd2;
        rom[190][19] = -8'd5;
        rom[190][20] = -8'd26;
        rom[190][21] = -8'd28;
        rom[190][22] = 8'd14;
        rom[190][23] = -8'd21;
        rom[190][24] = 8'd44;
        rom[190][25] = -8'd2;
        rom[190][26] = -8'd3;
        rom[190][27] = -8'd75;
        rom[190][28] = -8'd14;
        rom[190][29] = 8'd3;
        rom[190][30] = -8'd32;
        rom[190][31] = -8'd18;
        rom[191][0] = 8'd10;
        rom[191][1] = -8'd35;
        rom[191][2] = -8'd8;
        rom[191][3] = 8'd22;
        rom[191][4] = 8'd29;
        rom[191][5] = 8'd29;
        rom[191][6] = 8'd24;
        rom[191][7] = -8'd10;
        rom[191][8] = 8'd20;
        rom[191][9] = -8'd29;
        rom[191][10] = -8'd45;
        rom[191][11] = 8'd1;
        rom[191][12] = 8'd39;
        rom[191][13] = -8'd3;
        rom[191][14] = -8'd11;
        rom[191][15] = -8'd4;
        rom[191][16] = -8'd16;
        rom[191][17] = -8'd25;
        rom[191][18] = 8'd16;
        rom[191][19] = -8'd33;
        rom[191][20] = -8'd7;
        rom[191][21] = -8'd23;
        rom[191][22] = 8'd14;
        rom[191][23] = 8'd25;
        rom[191][24] = -8'd7;
        rom[191][25] = -8'd68;
        rom[191][26] = -8'd34;
        rom[191][27] = 8'd18;
        rom[191][28] = -8'd47;
        rom[191][29] = 8'd0;
        rom[191][30] = 8'd22;
        rom[191][31] = -8'd4;
        rom[192][0] = -8'd40;
        rom[192][1] = 8'd50;
        rom[192][2] = 8'd6;
        rom[192][3] = 8'd32;
        rom[192][4] = 8'd3;
        rom[192][5] = -8'd16;
        rom[192][6] = -8'd30;
        rom[192][7] = -8'd25;
        rom[192][8] = 8'd8;
        rom[192][9] = 8'd5;
        rom[192][10] = -8'd3;
        rom[192][11] = -8'd9;
        rom[192][12] = -8'd55;
        rom[192][13] = 8'd15;
        rom[192][14] = 8'd29;
        rom[192][15] = 8'd9;
        rom[192][16] = 8'd60;
        rom[192][17] = 8'd23;
        rom[192][18] = 8'd23;
        rom[192][19] = -8'd12;
        rom[192][20] = 8'd48;
        rom[192][21] = 8'd48;
        rom[192][22] = 8'd26;
        rom[192][23] = -8'd12;
        rom[192][24] = -8'd33;
        rom[192][25] = -8'd10;
        rom[192][26] = -8'd36;
        rom[192][27] = 8'd10;
        rom[192][28] = -8'd2;
        rom[192][29] = 8'd11;
        rom[192][30] = -8'd21;
        rom[192][31] = 8'd3;
        rom[193][0] = 8'd8;
        rom[193][1] = -8'd16;
        rom[193][2] = -8'd10;
        rom[193][3] = 8'd18;
        rom[193][4] = -8'd58;
        rom[193][5] = 8'd5;
        rom[193][6] = -8'd43;
        rom[193][7] = 8'd16;
        rom[193][8] = -8'd5;
        rom[193][9] = -8'd10;
        rom[193][10] = -8'd14;
        rom[193][11] = 8'd13;
        rom[193][12] = -8'd12;
        rom[193][13] = 8'd12;
        rom[193][14] = -8'd20;
        rom[193][15] = 8'd11;
        rom[193][16] = 8'd22;
        rom[193][17] = -8'd20;
        rom[193][18] = 8'd33;
        rom[193][19] = 8'd3;
        rom[193][20] = 8'd4;
        rom[193][21] = -8'd33;
        rom[193][22] = -8'd6;
        rom[193][23] = 8'd40;
        rom[193][24] = 8'd25;
        rom[193][25] = -8'd7;
        rom[193][26] = 8'd21;
        rom[193][27] = -8'd28;
        rom[193][28] = -8'd15;
        rom[193][29] = -8'd1;
        rom[193][30] = 8'd48;
        rom[193][31] = 8'd0;
        rom[194][0] = -8'd4;
        rom[194][1] = -8'd1;
        rom[194][2] = 8'd28;
        rom[194][3] = 8'd26;
        rom[194][4] = 8'd16;
        rom[194][5] = 8'd19;
        rom[194][6] = -8'd19;
        rom[194][7] = -8'd8;
        rom[194][8] = 8'd44;
        rom[194][9] = -8'd87;
        rom[194][10] = -8'd28;
        rom[194][11] = -8'd13;
        rom[194][12] = -8'd15;
        rom[194][13] = -8'd53;
        rom[194][14] = -8'd2;
        rom[194][15] = 8'd5;
        rom[194][16] = 8'd1;
        rom[194][17] = 8'd19;
        rom[194][18] = 8'd38;
        rom[194][19] = 8'd8;
        rom[194][20] = 8'd1;
        rom[194][21] = -8'd22;
        rom[194][22] = -8'd18;
        rom[194][23] = -8'd37;
        rom[194][24] = -8'd16;
        rom[194][25] = -8'd15;
        rom[194][26] = -8'd6;
        rom[194][27] = -8'd15;
        rom[194][28] = -8'd45;
        rom[194][29] = -8'd3;
        rom[194][30] = 8'd6;
        rom[194][31] = -8'd45;
        rom[195][0] = -8'd37;
        rom[195][1] = -8'd15;
        rom[195][2] = -8'd17;
        rom[195][3] = -8'd26;
        rom[195][4] = -8'd71;
        rom[195][5] = -8'd4;
        rom[195][6] = 8'd3;
        rom[195][7] = 8'd7;
        rom[195][8] = 8'd49;
        rom[195][9] = 8'd7;
        rom[195][10] = 8'd24;
        rom[195][11] = -8'd26;
        rom[195][12] = -8'd24;
        rom[195][13] = 8'd41;
        rom[195][14] = -8'd31;
        rom[195][15] = -8'd35;
        rom[195][16] = 8'd10;
        rom[195][17] = -8'd10;
        rom[195][18] = 8'd1;
        rom[195][19] = -8'd3;
        rom[195][20] = -8'd23;
        rom[195][21] = -8'd26;
        rom[195][22] = -8'd11;
        rom[195][23] = -8'd25;
        rom[195][24] = -8'd37;
        rom[195][25] = -8'd30;
        rom[195][26] = 8'd20;
        rom[195][27] = -8'd19;
        rom[195][28] = -8'd32;
        rom[195][29] = 8'd5;
        rom[195][30] = 8'd16;
        rom[195][31] = 8'd8;
        rom[196][0] = -8'd4;
        rom[196][1] = 8'd31;
        rom[196][2] = -8'd27;
        rom[196][3] = 8'd24;
        rom[196][4] = -8'd14;
        rom[196][5] = 8'd5;
        rom[196][6] = -8'd26;
        rom[196][7] = 8'd28;
        rom[196][8] = 8'd8;
        rom[196][9] = -8'd3;
        rom[196][10] = -8'd8;
        rom[196][11] = -8'd9;
        rom[196][12] = 8'd9;
        rom[196][13] = 8'd3;
        rom[196][14] = -8'd7;
        rom[196][15] = 8'd10;
        rom[196][16] = -8'd3;
        rom[196][17] = 8'd36;
        rom[196][18] = 8'd10;
        rom[196][19] = -8'd10;
        rom[196][20] = -8'd1;
        rom[196][21] = 8'd1;
        rom[196][22] = -8'd18;
        rom[196][23] = 8'd7;
        rom[196][24] = -8'd2;
        rom[196][25] = -8'd8;
        rom[196][26] = -8'd23;
        rom[196][27] = -8'd35;
        rom[196][28] = 8'd34;
        rom[196][29] = -8'd3;
        rom[196][30] = 8'd38;
        rom[196][31] = 8'd15;
        rom[197][0] = -8'd65;
        rom[197][1] = 8'd4;
        rom[197][2] = 8'd72;
        rom[197][3] = 8'd48;
        rom[197][4] = 8'd29;
        rom[197][5] = 8'd2;
        rom[197][6] = 8'd11;
        rom[197][7] = -8'd8;
        rom[197][8] = 8'd17;
        rom[197][9] = -8'd32;
        rom[197][10] = -8'd3;
        rom[197][11] = -8'd67;
        rom[197][12] = 8'd3;
        rom[197][13] = 8'd13;
        rom[197][14] = 8'd42;
        rom[197][15] = 8'd10;
        rom[197][16] = -8'd25;
        rom[197][17] = 8'd13;
        rom[197][18] = 8'd36;
        rom[197][19] = 8'd15;
        rom[197][20] = -8'd12;
        rom[197][21] = -8'd13;
        rom[197][22] = -8'd7;
        rom[197][23] = 8'd21;
        rom[197][24] = -8'd8;
        rom[197][25] = 8'd25;
        rom[197][26] = -8'd25;
        rom[197][27] = -8'd23;
        rom[197][28] = -8'd3;
        rom[197][29] = -8'd6;
        rom[197][30] = -8'd42;
        rom[197][31] = -8'd56;
        rom[198][0] = -8'd4;
        rom[198][1] = 8'd6;
        rom[198][2] = 8'd14;
        rom[198][3] = 8'd8;
        rom[198][4] = -8'd40;
        rom[198][5] = -8'd9;
        rom[198][6] = -8'd17;
        rom[198][7] = 8'd2;
        rom[198][8] = 8'd22;
        rom[198][9] = -8'd2;
        rom[198][10] = 8'd6;
        rom[198][11] = 8'd26;
        rom[198][12] = -8'd34;
        rom[198][13] = -8'd6;
        rom[198][14] = -8'd47;
        rom[198][15] = 8'd12;
        rom[198][16] = -8'd13;
        rom[198][17] = 8'd13;
        rom[198][18] = 8'd21;
        rom[198][19] = 8'd25;
        rom[198][20] = -8'd2;
        rom[198][21] = -8'd44;
        rom[198][22] = 8'd31;
        rom[198][23] = 8'd6;
        rom[198][24] = 8'd27;
        rom[198][25] = -8'd4;
        rom[198][26] = 8'd11;
        rom[198][27] = 8'd13;
        rom[198][28] = -8'd8;
        rom[198][29] = -8'd1;
        rom[198][30] = -8'd33;
        rom[198][31] = 8'd18;
        rom[199][0] = -8'd1;
        rom[199][1] = 8'd38;
        rom[199][2] = -8'd22;
        rom[199][3] = -8'd6;
        rom[199][4] = 8'd1;
        rom[199][5] = 8'd10;
        rom[199][6] = -8'd29;
        rom[199][7] = 8'd14;
        rom[199][8] = -8'd28;
        rom[199][9] = 8'd7;
        rom[199][10] = 8'd20;
        rom[199][11] = 8'd7;
        rom[199][12] = -8'd9;
        rom[199][13] = 8'd0;
        rom[199][14] = -8'd45;
        rom[199][15] = 8'd17;
        rom[199][16] = 8'd24;
        rom[199][17] = -8'd12;
        rom[199][18] = -8'd16;
        rom[199][19] = -8'd4;
        rom[199][20] = 8'd14;
        rom[199][21] = 8'd22;
        rom[199][22] = 8'd11;
        rom[199][23] = 8'd16;
        rom[199][24] = -8'd22;
        rom[199][25] = 8'd16;
        rom[199][26] = 8'd15;
        rom[199][27] = 8'd15;
        rom[199][28] = -8'd5;
        rom[199][29] = -8'd11;
        rom[199][30] = -8'd5;
        rom[199][31] = 8'd40;
        rom[200][0] = 8'd13;
        rom[200][1] = 8'd24;
        rom[200][2] = -8'd12;
        rom[200][3] = 8'd19;
        rom[200][4] = 8'd1;
        rom[200][5] = -8'd7;
        rom[200][6] = -8'd87;
        rom[200][7] = 8'd19;
        rom[200][8] = -8'd28;
        rom[200][9] = 8'd23;
        rom[200][10] = -8'd5;
        rom[200][11] = 8'd14;
        rom[200][12] = -8'd32;
        rom[200][13] = -8'd26;
        rom[200][14] = -8'd35;
        rom[200][15] = -8'd9;
        rom[200][16] = 8'd8;
        rom[200][17] = -8'd36;
        rom[200][18] = -8'd22;
        rom[200][19] = -8'd3;
        rom[200][20] = 8'd24;
        rom[200][21] = 8'd16;
        rom[200][22] = 8'd12;
        rom[200][23] = -8'd5;
        rom[200][24] = -8'd22;
        rom[200][25] = 8'd4;
        rom[200][26] = -8'd6;
        rom[200][27] = -8'd5;
        rom[200][28] = -8'd3;
        rom[200][29] = -8'd3;
        rom[200][30] = -8'd5;
        rom[200][31] = 8'd26;
        rom[201][0] = 8'd36;
        rom[201][1] = 8'd26;
        rom[201][2] = -8'd6;
        rom[201][3] = 8'd23;
        rom[201][4] = -8'd5;
        rom[201][5] = 8'd1;
        rom[201][6] = -8'd11;
        rom[201][7] = 8'd1;
        rom[201][8] = 8'd27;
        rom[201][9] = -8'd55;
        rom[201][10] = -8'd23;
        rom[201][11] = 8'd20;
        rom[201][12] = 8'd16;
        rom[201][13] = -8'd47;
        rom[201][14] = 8'd24;
        rom[201][15] = 8'd14;
        rom[201][16] = -8'd9;
        rom[201][17] = 8'd24;
        rom[201][18] = 8'd23;
        rom[201][19] = -8'd28;
        rom[201][20] = -8'd11;
        rom[201][21] = 8'd15;
        rom[201][22] = 8'd5;
        rom[201][23] = -8'd17;
        rom[201][24] = 8'd21;
        rom[201][25] = 8'd0;
        rom[201][26] = -8'd3;
        rom[201][27] = -8'd14;
        rom[201][28] = 8'd31;
        rom[201][29] = 8'd11;
        rom[201][30] = 8'd20;
        rom[201][31] = 8'd10;
        rom[202][0] = -8'd43;
        rom[202][1] = 8'd12;
        rom[202][2] = 8'd3;
        rom[202][3] = -8'd17;
        rom[202][4] = -8'd27;
        rom[202][5] = -8'd8;
        rom[202][6] = 8'd15;
        rom[202][7] = 8'd36;
        rom[202][8] = -8'd10;
        rom[202][9] = -8'd23;
        rom[202][10] = -8'd5;
        rom[202][11] = 8'd29;
        rom[202][12] = -8'd18;
        rom[202][13] = -8'd57;
        rom[202][14] = 8'd47;
        rom[202][15] = -8'd24;
        rom[202][16] = 8'd12;
        rom[202][17] = 8'd38;
        rom[202][18] = 8'd33;
        rom[202][19] = -8'd15;
        rom[202][20] = 8'd5;
        rom[202][21] = 8'd32;
        rom[202][22] = 8'd22;
        rom[202][23] = -8'd14;
        rom[202][24] = 8'd23;
        rom[202][25] = -8'd20;
        rom[202][26] = -8'd25;
        rom[202][27] = -8'd27;
        rom[202][28] = 8'd4;
        rom[202][29] = 8'd7;
        rom[202][30] = -8'd5;
        rom[202][31] = -8'd3;
        rom[203][0] = 8'd14;
        rom[203][1] = -8'd14;
        rom[203][2] = -8'd3;
        rom[203][3] = 8'd21;
        rom[203][4] = -8'd17;
        rom[203][5] = 8'd8;
        rom[203][6] = 8'd29;
        rom[203][7] = 8'd10;
        rom[203][8] = -8'd22;
        rom[203][9] = 8'd19;
        rom[203][10] = 8'd23;
        rom[203][11] = 8'd48;
        rom[203][12] = 8'd26;
        rom[203][13] = -8'd13;
        rom[203][14] = -8'd12;
        rom[203][15] = -8'd10;
        rom[203][16] = -8'd39;
        rom[203][17] = 8'd9;
        rom[203][18] = -8'd4;
        rom[203][19] = -8'd10;
        rom[203][20] = -8'd38;
        rom[203][21] = -8'd11;
        rom[203][22] = 8'd3;
        rom[203][23] = 8'd43;
        rom[203][24] = -8'd3;
        rom[203][25] = 8'd21;
        rom[203][26] = 8'd1;
        rom[203][27] = -8'd1;
        rom[203][28] = 8'd1;
        rom[203][29] = -8'd3;
        rom[203][30] = 8'd32;
        rom[203][31] = 8'd21;
        rom[204][0] = -8'd47;
        rom[204][1] = -8'd19;
        rom[204][2] = 8'd10;
        rom[204][3] = 8'd9;
        rom[204][4] = 8'd1;
        rom[204][5] = 8'd10;
        rom[204][6] = -8'd3;
        rom[204][7] = 8'd8;
        rom[204][8] = 8'd16;
        rom[204][9] = -8'd5;
        rom[204][10] = -8'd5;
        rom[204][11] = -8'd4;
        rom[204][12] = 8'd16;
        rom[204][13] = 8'd10;
        rom[204][14] = 8'd38;
        rom[204][15] = 8'd28;
        rom[204][16] = -8'd19;
        rom[204][17] = -8'd7;
        rom[204][18] = 8'd34;
        rom[204][19] = 8'd39;
        rom[204][20] = 8'd24;
        rom[204][21] = -8'd5;
        rom[204][22] = -8'd11;
        rom[204][23] = 8'd9;
        rom[204][24] = -8'd23;
        rom[204][25] = -8'd41;
        rom[204][26] = -8'd18;
        rom[204][27] = 8'd12;
        rom[204][28] = -8'd6;
        rom[204][29] = -8'd9;
        rom[204][30] = 8'd43;
        rom[204][31] = -8'd23;
        rom[205][0] = -8'd11;
        rom[205][1] = -8'd28;
        rom[205][2] = -8'd3;
        rom[205][3] = -8'd26;
        rom[205][4] = -8'd49;
        rom[205][5] = 8'd11;
        rom[205][6] = 8'd30;
        rom[205][7] = -8'd25;
        rom[205][8] = 8'd17;
        rom[205][9] = -8'd30;
        rom[205][10] = 8'd0;
        rom[205][11] = -8'd22;
        rom[205][12] = 8'd25;
        rom[205][13] = -8'd36;
        rom[205][14] = -8'd5;
        rom[205][15] = 8'd22;
        rom[205][16] = 8'd11;
        rom[205][17] = -8'd33;
        rom[205][18] = -8'd30;
        rom[205][19] = 8'd26;
        rom[205][20] = -8'd8;
        rom[205][21] = -8'd38;
        rom[205][22] = -8'd19;
        rom[205][23] = -8'd72;
        rom[205][24] = 8'd0;
        rom[205][25] = -8'd24;
        rom[205][26] = -8'd21;
        rom[205][27] = -8'd26;
        rom[205][28] = 8'd14;
        rom[205][29] = -8'd7;
        rom[205][30] = 8'd21;
        rom[205][31] = 8'd12;
        rom[206][0] = 8'd0;
        rom[206][1] = 8'd12;
        rom[206][2] = -8'd27;
        rom[206][3] = 8'd17;
        rom[206][4] = 8'd7;
        rom[206][5] = -8'd5;
        rom[206][6] = -8'd31;
        rom[206][7] = -8'd20;
        rom[206][8] = 8'd15;
        rom[206][9] = -8'd5;
        rom[206][10] = -8'd29;
        rom[206][11] = -8'd15;
        rom[206][12] = -8'd2;
        rom[206][13] = 8'd3;
        rom[206][14] = -8'd24;
        rom[206][15] = 8'd22;
        rom[206][16] = 8'd1;
        rom[206][17] = -8'd15;
        rom[206][18] = -8'd13;
        rom[206][19] = -8'd3;
        rom[206][20] = 8'd18;
        rom[206][21] = 8'd4;
        rom[206][22] = -8'd23;
        rom[206][23] = -8'd2;
        rom[206][24] = -8'd28;
        rom[206][25] = 8'd10;
        rom[206][26] = 8'd1;
        rom[206][27] = 8'd1;
        rom[206][28] = 8'd6;
        rom[206][29] = 8'd1;
        rom[206][30] = 8'd23;
        rom[206][31] = 8'd33;
        rom[207][0] = -8'd59;
        rom[207][1] = 8'd61;
        rom[207][2] = -8'd18;
        rom[207][3] = 8'd3;
        rom[207][4] = -8'd7;
        rom[207][5] = -8'd24;
        rom[207][6] = 8'd5;
        rom[207][7] = -8'd45;
        rom[207][8] = 8'd31;
        rom[207][9] = -8'd20;
        rom[207][10] = -8'd7;
        rom[207][11] = -8'd32;
        rom[207][12] = -8'd45;
        rom[207][13] = -8'd2;
        rom[207][14] = 8'd18;
        rom[207][15] = 8'd28;
        rom[207][16] = 8'd38;
        rom[207][17] = -8'd29;
        rom[207][18] = -8'd19;
        rom[207][19] = -8'd7;
        rom[207][20] = -8'd7;
        rom[207][21] = 8'd35;
        rom[207][22] = 8'd10;
        rom[207][23] = -8'd29;
        rom[207][24] = -8'd49;
        rom[207][25] = 8'd26;
        rom[207][26] = 8'd25;
        rom[207][27] = 8'd11;
        rom[207][28] = -8'd11;
        rom[207][29] = -8'd9;
        rom[207][30] = -8'd9;
        rom[207][31] = 8'd3;
        rom[208][0] = -8'd4;
        rom[208][1] = 8'd22;
        rom[208][2] = 8'd0;
        rom[208][3] = -8'd15;
        rom[208][4] = -8'd16;
        rom[208][5] = 8'd5;
        rom[208][6] = -8'd24;
        rom[208][7] = 8'd1;
        rom[208][8] = 8'd3;
        rom[208][9] = 8'd7;
        rom[208][10] = 8'd37;
        rom[208][11] = 8'd2;
        rom[208][12] = -8'd16;
        rom[208][13] = 8'd3;
        rom[208][14] = 8'd25;
        rom[208][15] = -8'd16;
        rom[208][16] = 8'd4;
        rom[208][17] = 8'd8;
        rom[208][18] = 8'd3;
        rom[208][19] = -8'd89;
        rom[208][20] = -8'd24;
        rom[208][21] = -8'd25;
        rom[208][22] = -8'd4;
        rom[208][23] = -8'd25;
        rom[208][24] = -8'd37;
        rom[208][25] = -8'd61;
        rom[208][26] = 8'd1;
        rom[208][27] = -8'd12;
        rom[208][28] = -8'd4;
        rom[208][29] = -8'd8;
        rom[208][30] = -8'd3;
        rom[208][31] = 8'd11;
        rom[209][0] = -8'd8;
        rom[209][1] = -8'd13;
        rom[209][2] = 8'd1;
        rom[209][3] = -8'd41;
        rom[209][4] = -8'd4;
        rom[209][5] = -8'd4;
        rom[209][6] = -8'd31;
        rom[209][7] = -8'd13;
        rom[209][8] = 8'd12;
        rom[209][9] = -8'd23;
        rom[209][10] = 8'd5;
        rom[209][11] = -8'd27;
        rom[209][12] = -8'd35;
        rom[209][13] = -8'd60;
        rom[209][14] = 8'd14;
        rom[209][15] = -8'd13;
        rom[209][16] = 8'd27;
        rom[209][17] = 8'd25;
        rom[209][18] = -8'd17;
        rom[209][19] = 8'd12;
        rom[209][20] = 8'd25;
        rom[209][21] = -8'd4;
        rom[209][22] = 8'd15;
        rom[209][23] = -8'd23;
        rom[209][24] = -8'd18;
        rom[209][25] = -8'd13;
        rom[209][26] = -8'd19;
        rom[209][27] = 8'd1;
        rom[209][28] = -8'd26;
        rom[209][29] = -8'd8;
        rom[209][30] = -8'd23;
        rom[209][31] = -8'd24;
        rom[210][0] = -8'd24;
        rom[210][1] = 8'd28;
        rom[210][2] = 8'd7;
        rom[210][3] = 8'd2;
        rom[210][4] = -8'd34;
        rom[210][5] = -8'd11;
        rom[210][6] = 8'd4;
        rom[210][7] = -8'd8;
        rom[210][8] = 8'd9;
        rom[210][9] = -8'd9;
        rom[210][10] = -8'd17;
        rom[210][11] = -8'd31;
        rom[210][12] = -8'd5;
        rom[210][13] = -8'd2;
        rom[210][14] = 8'd12;
        rom[210][15] = 8'd34;
        rom[210][16] = 8'd41;
        rom[210][17] = -8'd30;
        rom[210][18] = 8'd21;
        rom[210][19] = 8'd26;
        rom[210][20] = 8'd6;
        rom[210][21] = 8'd35;
        rom[210][22] = -8'd34;
        rom[210][23] = -8'd35;
        rom[210][24] = -8'd35;
        rom[210][25] = -8'd10;
        rom[210][26] = -8'd3;
        rom[210][27] = 8'd12;
        rom[210][28] = 8'd35;
        rom[210][29] = 8'd5;
        rom[210][30] = -8'd9;
        rom[210][31] = 8'd34;
        rom[211][0] = -8'd52;
        rom[211][1] = 8'd2;
        rom[211][2] = -8'd40;
        rom[211][3] = 8'd29;
        rom[211][4] = -8'd26;
        rom[211][5] = 8'd7;
        rom[211][6] = -8'd16;
        rom[211][7] = -8'd12;
        rom[211][8] = 8'd8;
        rom[211][9] = -8'd3;
        rom[211][10] = -8'd16;
        rom[211][11] = -8'd15;
        rom[211][12] = 8'd37;
        rom[211][13] = 8'd6;
        rom[211][14] = 8'd6;
        rom[211][15] = 8'd12;
        rom[211][16] = -8'd31;
        rom[211][17] = -8'd6;
        rom[211][18] = 8'd4;
        rom[211][19] = -8'd2;
        rom[211][20] = 8'd3;
        rom[211][21] = 8'd17;
        rom[211][22] = -8'd3;
        rom[211][23] = -8'd7;
        rom[211][24] = -8'd10;
        rom[211][25] = 8'd22;
        rom[211][26] = 8'd9;
        rom[211][27] = -8'd33;
        rom[211][28] = -8'd1;
        rom[211][29] = -8'd9;
        rom[211][30] = -8'd16;
        rom[211][31] = -8'd40;
        rom[212][0] = 8'd13;
        rom[212][1] = 8'd1;
        rom[212][2] = -8'd2;
        rom[212][3] = -8'd2;
        rom[212][4] = 8'd57;
        rom[212][5] = -8'd2;
        rom[212][6] = -8'd48;
        rom[212][7] = -8'd31;
        rom[212][8] = 8'd8;
        rom[212][9] = -8'd8;
        rom[212][10] = 8'd10;
        rom[212][11] = 8'd9;
        rom[212][12] = 8'd30;
        rom[212][13] = -8'd19;
        rom[212][14] = -8'd32;
        rom[212][15] = -8'd19;
        rom[212][16] = -8'd31;
        rom[212][17] = 8'd5;
        rom[212][18] = -8'd9;
        rom[212][19] = -8'd45;
        rom[212][20] = -8'd26;
        rom[212][21] = 8'd19;
        rom[212][22] = 8'd3;
        rom[212][23] = 8'd30;
        rom[212][24] = -8'd1;
        rom[212][25] = -8'd7;
        rom[212][26] = -8'd23;
        rom[212][27] = -8'd6;
        rom[212][28] = -8'd24;
        rom[212][29] = 8'd2;
        rom[212][30] = -8'd13;
        rom[212][31] = -8'd38;
        rom[213][0] = 8'd38;
        rom[213][1] = -8'd17;
        rom[213][2] = -8'd15;
        rom[213][3] = 8'd21;
        rom[213][4] = 8'd48;
        rom[213][5] = 8'd41;
        rom[213][6] = 8'd13;
        rom[213][7] = -8'd25;
        rom[213][8] = 8'd14;
        rom[213][9] = 8'd20;
        rom[213][10] = -8'd10;
        rom[213][11] = -8'd1;
        rom[213][12] = -8'd12;
        rom[213][13] = 8'd5;
        rom[213][14] = -8'd4;
        rom[213][15] = -8'd14;
        rom[213][16] = -8'd46;
        rom[213][17] = -8'd19;
        rom[213][18] = -8'd8;
        rom[213][19] = 8'd9;
        rom[213][20] = -8'd16;
        rom[213][21] = -8'd1;
        rom[213][22] = 8'd22;
        rom[213][23] = 8'd17;
        rom[213][24] = 8'd34;
        rom[213][25] = 8'd17;
        rom[213][26] = -8'd21;
        rom[213][27] = -8'd6;
        rom[213][28] = -8'd17;
        rom[213][29] = 8'd4;
        rom[213][30] = 8'd16;
        rom[213][31] = 8'd4;
        rom[214][0] = -8'd26;
        rom[214][1] = -8'd18;
        rom[214][2] = -8'd12;
        rom[214][3] = 8'd31;
        rom[214][4] = 8'd23;
        rom[214][5] = -8'd32;
        rom[214][6] = -8'd12;
        rom[214][7] = 8'd5;
        rom[214][8] = 8'd6;
        rom[214][9] = 8'd9;
        rom[214][10] = 8'd2;
        rom[214][11] = -8'd11;
        rom[214][12] = -8'd25;
        rom[214][13] = -8'd11;
        rom[214][14] = 8'd16;
        rom[214][15] = -8'd19;
        rom[214][16] = 8'd25;
        rom[214][17] = 8'd30;
        rom[214][18] = 8'd6;
        rom[214][19] = 8'd34;
        rom[214][20] = -8'd11;
        rom[214][21] = -8'd3;
        rom[214][22] = 8'd21;
        rom[214][23] = -8'd16;
        rom[214][24] = -8'd44;
        rom[214][25] = -8'd43;
        rom[214][26] = 8'd1;
        rom[214][27] = -8'd16;
        rom[214][28] = -8'd23;
        rom[214][29] = -8'd10;
        rom[214][30] = 8'd7;
        rom[214][31] = -8'd3;
        rom[215][0] = 8'd5;
        rom[215][1] = -8'd38;
        rom[215][2] = 8'd16;
        rom[215][3] = 8'd11;
        rom[215][4] = -8'd13;
        rom[215][5] = -8'd17;
        rom[215][6] = -8'd36;
        rom[215][7] = -8'd1;
        rom[215][8] = -8'd24;
        rom[215][9] = 8'd15;
        rom[215][10] = -8'd12;
        rom[215][11] = -8'd17;
        rom[215][12] = -8'd20;
        rom[215][13] = -8'd23;
        rom[215][14] = 8'd32;
        rom[215][15] = -8'd19;
        rom[215][16] = 8'd9;
        rom[215][17] = -8'd8;
        rom[215][18] = 8'd2;
        rom[215][19] = -8'd2;
        rom[215][20] = 8'd1;
        rom[215][21] = -8'd33;
        rom[215][22] = -8'd74;
        rom[215][23] = 8'd11;
        rom[215][24] = -8'd3;
        rom[215][25] = -8'd19;
        rom[215][26] = -8'd4;
        rom[215][27] = -8'd30;
        rom[215][28] = -8'd3;
        rom[215][29] = 8'd1;
        rom[215][30] = -8'd2;
        rom[215][31] = 8'd29;
        rom[216][0] = 8'd40;
        rom[216][1] = 8'd6;
        rom[216][2] = 8'd36;
        rom[216][3] = 8'd33;
        rom[216][4] = -8'd14;
        rom[216][5] = 8'd19;
        rom[216][6] = 8'd13;
        rom[216][7] = 8'd16;
        rom[216][8] = 8'd4;
        rom[216][9] = -8'd11;
        rom[216][10] = -8'd33;
        rom[216][11] = -8'd68;
        rom[216][12] = 8'd10;
        rom[216][13] = 8'd55;
        rom[216][14] = 8'd12;
        rom[216][15] = 8'd19;
        rom[216][16] = -8'd40;
        rom[216][17] = -8'd49;
        rom[216][18] = -8'd3;
        rom[216][19] = -8'd24;
        rom[216][20] = 8'd31;
        rom[216][21] = 8'd28;
        rom[216][22] = -8'd97;
        rom[216][23] = 8'd10;
        rom[216][24] = 8'd3;
        rom[216][25] = 8'd24;
        rom[216][26] = -8'd36;
        rom[216][27] = 8'd1;
        rom[216][28] = -8'd6;
        rom[216][29] = -8'd10;
        rom[216][30] = -8'd3;
        rom[216][31] = -8'd18;
        rom[217][0] = 8'd35;
        rom[217][1] = 8'd4;
        rom[217][2] = -8'd6;
        rom[217][3] = 8'd12;
        rom[217][4] = 8'd7;
        rom[217][5] = -8'd12;
        rom[217][6] = -8'd12;
        rom[217][7] = 8'd18;
        rom[217][8] = 8'd4;
        rom[217][9] = 8'd11;
        rom[217][10] = 8'd11;
        rom[217][11] = -8'd57;
        rom[217][12] = -8'd6;
        rom[217][13] = 8'd8;
        rom[217][14] = 8'd28;
        rom[217][15] = 8'd4;
        rom[217][16] = 8'd38;
        rom[217][17] = 8'd14;
        rom[217][18] = -8'd20;
        rom[217][19] = -8'd1;
        rom[217][20] = 8'd2;
        rom[217][21] = 8'd30;
        rom[217][22] = 8'd14;
        rom[217][23] = 8'd2;
        rom[217][24] = 8'd5;
        rom[217][25] = -8'd42;
        rom[217][26] = 8'd1;
        rom[217][27] = 8'd19;
        rom[217][28] = 8'd12;
        rom[217][29] = -8'd3;
        rom[217][30] = -8'd34;
        rom[217][31] = -8'd9;
        rom[218][0] = 8'd2;
        rom[218][1] = -8'd32;
        rom[218][2] = 8'd30;
        rom[218][3] = 8'd20;
        rom[218][4] = 8'd8;
        rom[218][5] = 8'd16;
        rom[218][6] = 8'd32;
        rom[218][7] = 8'd3;
        rom[218][8] = -8'd7;
        rom[218][9] = 8'd21;
        rom[218][10] = -8'd13;
        rom[218][11] = -8'd2;
        rom[218][12] = 8'd3;
        rom[218][13] = -8'd28;
        rom[218][14] = -8'd21;
        rom[218][15] = 8'd22;
        rom[218][16] = 8'd20;
        rom[218][17] = 8'd1;
        rom[218][18] = 8'd12;
        rom[218][19] = 8'd10;
        rom[218][20] = 8'd10;
        rom[218][21] = 8'd17;
        rom[218][22] = -8'd4;
        rom[218][23] = 8'd7;
        rom[218][24] = -8'd22;
        rom[218][25] = -8'd11;
        rom[218][26] = -8'd9;
        rom[218][27] = -8'd16;
        rom[218][28] = 8'd3;
        rom[218][29] = -8'd5;
        rom[218][30] = 8'd12;
        rom[218][31] = 8'd2;
        rom[219][0] = 8'd19;
        rom[219][1] = 8'd19;
        rom[219][2] = -8'd16;
        rom[219][3] = -8'd12;
        rom[219][4] = -8'd33;
        rom[219][5] = 8'd9;
        rom[219][6] = -8'd18;
        rom[219][7] = 8'd0;
        rom[219][8] = -8'd9;
        rom[219][9] = -8'd4;
        rom[219][10] = 8'd2;
        rom[219][11] = 8'd25;
        rom[219][12] = 8'd1;
        rom[219][13] = 8'd13;
        rom[219][14] = -8'd6;
        rom[219][15] = 8'd21;
        rom[219][16] = -8'd7;
        rom[219][17] = -8'd23;
        rom[219][18] = -8'd1;
        rom[219][19] = -8'd17;
        rom[219][20] = 8'd42;
        rom[219][21] = 8'd17;
        rom[219][22] = -8'd7;
        rom[219][23] = 8'd4;
        rom[219][24] = -8'd18;
        rom[219][25] = 8'd32;
        rom[219][26] = 8'd16;
        rom[219][27] = -8'd8;
        rom[219][28] = 8'd13;
        rom[219][29] = 8'd3;
        rom[219][30] = 8'd31;
        rom[219][31] = 8'd40;
        rom[220][0] = -8'd19;
        rom[220][1] = -8'd1;
        rom[220][2] = -8'd2;
        rom[220][3] = -8'd9;
        rom[220][4] = -8'd1;
        rom[220][5] = 8'd10;
        rom[220][6] = 8'd15;
        rom[220][7] = 8'd10;
        rom[220][8] = 8'd22;
        rom[220][9] = -8'd13;
        rom[220][10] = -8'd4;
        rom[220][11] = -8'd1;
        rom[220][12] = -8'd57;
        rom[220][13] = -8'd46;
        rom[220][14] = 8'd29;
        rom[220][15] = -8'd29;
        rom[220][16] = -8'd6;
        rom[220][17] = -8'd3;
        rom[220][18] = 8'd28;
        rom[220][19] = -8'd11;
        rom[220][20] = -8'd40;
        rom[220][21] = 8'd22;
        rom[220][22] = 8'd15;
        rom[220][23] = -8'd47;
        rom[220][24] = -8'd17;
        rom[220][25] = -8'd11;
        rom[220][26] = -8'd25;
        rom[220][27] = 8'd25;
        rom[220][28] = -8'd12;
        rom[220][29] = -8'd1;
        rom[220][30] = -8'd20;
        rom[220][31] = -8'd71;
        rom[221][0] = 8'd25;
        rom[221][1] = -8'd16;
        rom[221][2] = -8'd2;
        rom[221][3] = -8'd1;
        rom[221][4] = 8'd19;
        rom[221][5] = -8'd47;
        rom[221][6] = 8'd13;
        rom[221][7] = -8'd42;
        rom[221][8] = -8'd23;
        rom[221][9] = -8'd25;
        rom[221][10] = -8'd19;
        rom[221][11] = -8'd18;
        rom[221][12] = 8'd38;
        rom[221][13] = -8'd7;
        rom[221][14] = -8'd18;
        rom[221][15] = 8'd1;
        rom[221][16] = -8'd15;
        rom[221][17] = 8'd14;
        rom[221][18] = 8'd45;
        rom[221][19] = 8'd5;
        rom[221][20] = 8'd8;
        rom[221][21] = -8'd29;
        rom[221][22] = -8'd2;
        rom[221][23] = 8'd11;
        rom[221][24] = 8'd14;
        rom[221][25] = 8'd13;
        rom[221][26] = 8'd1;
        rom[221][27] = -8'd9;
        rom[221][28] = -8'd18;
        rom[221][29] = -8'd12;
        rom[221][30] = 8'd2;
        rom[221][31] = -8'd7;
        rom[222][0] = 8'd7;
        rom[222][1] = 8'd38;
        rom[222][2] = 8'd29;
        rom[222][3] = 8'd3;
        rom[222][4] = 8'd27;
        rom[222][5] = 8'd17;
        rom[222][6] = 8'd9;
        rom[222][7] = 8'd16;
        rom[222][8] = -8'd14;
        rom[222][9] = 8'd23;
        rom[222][10] = 8'd16;
        rom[222][11] = 8'd30;
        rom[222][12] = -8'd57;
        rom[222][13] = 8'd0;
        rom[222][14] = 8'd15;
        rom[222][15] = 8'd34;
        rom[222][16] = -8'd4;
        rom[222][17] = 8'd18;
        rom[222][18] = 8'd20;
        rom[222][19] = -8'd17;
        rom[222][20] = 8'd6;
        rom[222][21] = 8'd64;
        rom[222][22] = 8'd26;
        rom[222][23] = -8'd26;
        rom[222][24] = -8'd19;
        rom[222][25] = 8'd5;
        rom[222][26] = -8'd21;
        rom[222][27] = 8'd35;
        rom[222][28] = 8'd33;
        rom[222][29] = 8'd10;
        rom[222][30] = 8'd6;
        rom[222][31] = -8'd38;
        rom[223][0] = 8'd10;
        rom[223][1] = 8'd35;
        rom[223][2] = 8'd33;
        rom[223][3] = -8'd19;
        rom[223][4] = 8'd9;
        rom[223][5] = 8'd26;
        rom[223][6] = -8'd41;
        rom[223][7] = 8'd6;
        rom[223][8] = -8'd29;
        rom[223][9] = -8'd45;
        rom[223][10] = -8'd44;
        rom[223][11] = -8'd20;
        rom[223][12] = 8'd17;
        rom[223][13] = -8'd27;
        rom[223][14] = -8'd40;
        rom[223][15] = -8'd18;
        rom[223][16] = -8'd25;
        rom[223][17] = -8'd44;
        rom[223][18] = -8'd22;
        rom[223][19] = 8'd19;
        rom[223][20] = -8'd38;
        rom[223][21] = 8'd60;
        rom[223][22] = -8'd53;
        rom[223][23] = -8'd58;
        rom[223][24] = -8'd25;
        rom[223][25] = 8'd59;
        rom[223][26] = 8'd16;
        rom[223][27] = -8'd26;
        rom[223][28] = -8'd12;
        rom[223][29] = 8'd4;
        rom[223][30] = -8'd48;
        rom[223][31] = -8'd24;
        rom[224][0] = -8'd37;
        rom[224][1] = -8'd12;
        rom[224][2] = 8'd8;
        rom[224][3] = -8'd4;
        rom[224][4] = -8'd38;
        rom[224][5] = 8'd25;
        rom[224][6] = -8'd24;
        rom[224][7] = -8'd26;
        rom[224][8] = 8'd6;
        rom[224][9] = 8'd13;
        rom[224][10] = 8'd10;
        rom[224][11] = 8'd15;
        rom[224][12] = -8'd65;
        rom[224][13] = 8'd10;
        rom[224][14] = 8'd38;
        rom[224][15] = -8'd32;
        rom[224][16] = 8'd35;
        rom[224][17] = -8'd9;
        rom[224][18] = 8'd9;
        rom[224][19] = -8'd15;
        rom[224][20] = 8'd9;
        rom[224][21] = -8'd14;
        rom[224][22] = 8'd36;
        rom[224][23] = -8'd9;
        rom[224][24] = -8'd25;
        rom[224][25] = 8'd2;
        rom[224][26] = -8'd48;
        rom[224][27] = 8'd32;
        rom[224][28] = 8'd3;
        rom[224][29] = -8'd3;
        rom[224][30] = 8'd2;
        rom[224][31] = -8'd3;
        rom[225][0] = -8'd11;
        rom[225][1] = 8'd20;
        rom[225][2] = -8'd21;
        rom[225][3] = 8'd2;
        rom[225][4] = -8'd56;
        rom[225][5] = 8'd26;
        rom[225][6] = -8'd37;
        rom[225][7] = 8'd28;
        rom[225][8] = -8'd2;
        rom[225][9] = 8'd23;
        rom[225][10] = -8'd4;
        rom[225][11] = 8'd1;
        rom[225][12] = 8'd4;
        rom[225][13] = -8'd30;
        rom[225][14] = -8'd4;
        rom[225][15] = 8'd4;
        rom[225][16] = 8'd39;
        rom[225][17] = -8'd16;
        rom[225][18] = -8'd4;
        rom[225][19] = 8'd7;
        rom[225][20] = 8'd33;
        rom[225][21] = 8'd22;
        rom[225][22] = 8'd18;
        rom[225][23] = 8'd10;
        rom[225][24] = 8'd11;
        rom[225][25] = -8'd29;
        rom[225][26] = -8'd6;
        rom[225][27] = -8'd24;
        rom[225][28] = -8'd28;
        rom[225][29] = -8'd2;
        rom[225][30] = 8'd17;
        rom[225][31] = 8'd41;
        rom[226][0] = -8'd2;
        rom[226][1] = -8'd5;
        rom[226][2] = 8'd8;
        rom[226][3] = 8'd49;
        rom[226][4] = -8'd14;
        rom[226][5] = 8'd4;
        rom[226][6] = 8'd3;
        rom[226][7] = 8'd8;
        rom[226][8] = -8'd20;
        rom[226][9] = -8'd62;
        rom[226][10] = -8'd29;
        rom[226][11] = 8'd2;
        rom[226][12] = 8'd14;
        rom[226][13] = -8'd62;
        rom[226][14] = -8'd14;
        rom[226][15] = -8'd11;
        rom[226][16] = -8'd25;
        rom[226][17] = 8'd34;
        rom[226][18] = 8'd10;
        rom[226][19] = -8'd1;
        rom[226][20] = -8'd37;
        rom[226][21] = -8'd12;
        rom[226][22] = -8'd10;
        rom[226][23] = 8'd15;
        rom[226][24] = 8'd2;
        rom[226][25] = 8'd7;
        rom[226][26] = 8'd14;
        rom[226][27] = -8'd34;
        rom[226][28] = -8'd20;
        rom[226][29] = 8'd4;
        rom[226][30] = 8'd21;
        rom[226][31] = -8'd4;
        rom[227][0] = -8'd3;
        rom[227][1] = -8'd45;
        rom[227][2] = 8'd17;
        rom[227][3] = -8'd10;
        rom[227][4] = -8'd70;
        rom[227][5] = -8'd12;
        rom[227][6] = -8'd10;
        rom[227][7] = -8'd8;
        rom[227][8] = 8'd2;
        rom[227][9] = -8'd12;
        rom[227][10] = -8'd14;
        rom[227][11] = 8'd12;
        rom[227][12] = -8'd58;
        rom[227][13] = 8'd23;
        rom[227][14] = -8'd40;
        rom[227][15] = -8'd38;
        rom[227][16] = -8'd37;
        rom[227][17] = 8'd6;
        rom[227][18] = 8'd4;
        rom[227][19] = -8'd30;
        rom[227][20] = -8'd11;
        rom[227][21] = -8'd58;
        rom[227][22] = 8'd20;
        rom[227][23] = -8'd2;
        rom[227][24] = 8'd12;
        rom[227][25] = -8'd41;
        rom[227][26] = 8'd23;
        rom[227][27] = -8'd9;
        rom[227][28] = -8'd34;
        rom[227][29] = -8'd8;
        rom[227][30] = 8'd30;
        rom[227][31] = -8'd26;
        rom[228][0] = -8'd21;
        rom[228][1] = 8'd1;
        rom[228][2] = 8'd2;
        rom[228][3] = -8'd28;
        rom[228][4] = -8'd27;
        rom[228][5] = 8'd12;
        rom[228][6] = -8'd27;
        rom[228][7] = 8'd50;
        rom[228][8] = 8'd11;
        rom[228][9] = 8'd5;
        rom[228][10] = 8'd6;
        rom[228][11] = 8'd28;
        rom[228][12] = 8'd12;
        rom[228][13] = -8'd9;
        rom[228][14] = 8'd38;
        rom[228][15] = 8'd38;
        rom[228][16] = 8'd11;
        rom[228][17] = 8'd6;
        rom[228][18] = -8'd26;
        rom[228][19] = -8'd35;
        rom[228][20] = 8'd18;
        rom[228][21] = 8'd21;
        rom[228][22] = 8'd36;
        rom[228][23] = -8'd47;
        rom[228][24] = -8'd2;
        rom[228][25] = -8'd33;
        rom[228][26] = -8'd29;
        rom[228][27] = -8'd1;
        rom[228][28] = -8'd22;
        rom[228][29] = 8'd4;
        rom[228][30] = 8'd46;
        rom[228][31] = 8'd6;
        rom[229][0] = -8'd39;
        rom[229][1] = 8'd3;
        rom[229][2] = 8'd33;
        rom[229][3] = 8'd0;
        rom[229][4] = 8'd59;
        rom[229][5] = -8'd5;
        rom[229][6] = 8'd3;
        rom[229][7] = -8'd33;
        rom[229][8] = -8'd51;
        rom[229][9] = -8'd22;
        rom[229][10] = -8'd22;
        rom[229][11] = -8'd44;
        rom[229][12] = -8'd41;
        rom[229][13] = 8'd8;
        rom[229][14] = 8'd19;
        rom[229][15] = -8'd81;
        rom[229][16] = 8'd30;
        rom[229][17] = 8'd45;
        rom[229][18] = -8'd36;
        rom[229][19] = 8'd6;
        rom[229][20] = -8'd27;
        rom[229][21] = 8'd17;
        rom[229][22] = -8'd13;
        rom[229][23] = 8'd37;
        rom[229][24] = 8'd30;
        rom[229][25] = -8'd13;
        rom[229][26] = -8'd30;
        rom[229][27] = -8'd52;
        rom[229][28] = -8'd9;
        rom[229][29] = -8'd1;
        rom[229][30] = -8'd56;
        rom[229][31] = -8'd33;
        rom[230][0] = 8'd8;
        rom[230][1] = -8'd10;
        rom[230][2] = 8'd22;
        rom[230][3] = -8'd10;
        rom[230][4] = -8'd16;
        rom[230][5] = 8'd31;
        rom[230][6] = -8'd21;
        rom[230][7] = -8'd14;
        rom[230][8] = 8'd15;
        rom[230][9] = -8'd19;
        rom[230][10] = -8'd21;
        rom[230][11] = -8'd12;
        rom[230][12] = -8'd55;
        rom[230][13] = 8'd26;
        rom[230][14] = -8'd23;
        rom[230][15] = -8'd2;
        rom[230][16] = 8'd23;
        rom[230][17] = -8'd5;
        rom[230][18] = -8'd8;
        rom[230][19] = 8'd32;
        rom[230][20] = 8'd2;
        rom[230][21] = -8'd51;
        rom[230][22] = 8'd22;
        rom[230][23] = -8'd9;
        rom[230][24] = 8'd3;
        rom[230][25] = -8'd25;
        rom[230][26] = 8'd16;
        rom[230][27] = -8'd1;
        rom[230][28] = 8'd28;
        rom[230][29] = 8'd7;
        rom[230][30] = -8'd8;
        rom[230][31] = -8'd15;
        rom[231][0] = 8'd19;
        rom[231][1] = 8'd30;
        rom[231][2] = -8'd34;
        rom[231][3] = -8'd3;
        rom[231][4] = -8'd18;
        rom[231][5] = -8'd24;
        rom[231][6] = -8'd31;
        rom[231][7] = 8'd5;
        rom[231][8] = 8'd17;
        rom[231][9] = 8'd1;
        rom[231][10] = 8'd23;
        rom[231][11] = 8'd11;
        rom[231][12] = 8'd9;
        rom[231][13] = 8'd23;
        rom[231][14] = -8'd78;
        rom[231][15] = 8'd7;
        rom[231][16] = 8'd0;
        rom[231][17] = -8'd19;
        rom[231][18] = 8'd13;
        rom[231][19] = -8'd2;
        rom[231][20] = -8'd1;
        rom[231][21] = 8'd0;
        rom[231][22] = 8'd24;
        rom[231][23] = -8'd23;
        rom[231][24] = -8'd4;
        rom[231][25] = 8'd17;
        rom[231][26] = 8'd19;
        rom[231][27] = 8'd4;
        rom[231][28] = -8'd7;
        rom[231][29] = -8'd5;
        rom[231][30] = -8'd14;
        rom[231][31] = 8'd34;
        rom[232][0] = 8'd0;
        rom[232][1] = 8'd5;
        rom[232][2] = 8'd2;
        rom[232][3] = 8'd6;
        rom[232][4] = -8'd27;
        rom[232][5] = -8'd15;
        rom[232][6] = -8'd61;
        rom[232][7] = 8'd11;
        rom[232][8] = -8'd11;
        rom[232][9] = 8'd7;
        rom[232][10] = 8'd13;
        rom[232][11] = 8'd22;
        rom[232][12] = -8'd39;
        rom[232][13] = -8'd30;
        rom[232][14] = -8'd18;
        rom[232][15] = -8'd22;
        rom[232][16] = -8'd29;
        rom[232][17] = 8'd39;
        rom[232][18] = -8'd26;
        rom[232][19] = -8'd15;
        rom[232][20] = -8'd10;
        rom[232][21] = -8'd6;
        rom[232][22] = -8'd19;
        rom[232][23] = -8'd29;
        rom[232][24] = -8'd22;
        rom[232][25] = -8'd19;
        rom[232][26] = 8'd1;
        rom[232][27] = -8'd7;
        rom[232][28] = -8'd40;
        rom[232][29] = -8'd14;
        rom[232][30] = -8'd30;
        rom[232][31] = 8'd12;
        rom[233][0] = 8'd15;
        rom[233][1] = -8'd20;
        rom[233][2] = -8'd38;
        rom[233][3] = 8'd19;
        rom[233][4] = -8'd17;
        rom[233][5] = 8'd33;
        rom[233][6] = -8'd23;
        rom[233][7] = -8'd38;
        rom[233][8] = -8'd36;
        rom[233][9] = -8'd26;
        rom[233][10] = -8'd56;
        rom[233][11] = 8'd34;
        rom[233][12] = -8'd9;
        rom[233][13] = -8'd6;
        rom[233][14] = -8'd29;
        rom[233][15] = -8'd7;
        rom[233][16] = -8'd24;
        rom[233][17] = -8'd45;
        rom[233][18] = -8'd3;
        rom[233][19] = -8'd33;
        rom[233][20] = -8'd25;
        rom[233][21] = -8'd31;
        rom[233][22] = 8'd0;
        rom[233][23] = 8'd48;
        rom[233][24] = 8'd23;
        rom[233][25] = -8'd24;
        rom[233][26] = -8'd20;
        rom[233][27] = -8'd1;
        rom[233][28] = 8'd31;
        rom[233][29] = 8'd1;
        rom[233][30] = 8'd19;
        rom[233][31] = 8'd35;
        rom[234][0] = -8'd41;
        rom[234][1] = -8'd5;
        rom[234][2] = -8'd19;
        rom[234][3] = 8'd16;
        rom[234][4] = -8'd22;
        rom[234][5] = -8'd2;
        rom[234][6] = -8'd55;
        rom[234][7] = 8'd24;
        rom[234][8] = 8'd15;
        rom[234][9] = -8'd23;
        rom[234][10] = -8'd4;
        rom[234][11] = 8'd60;
        rom[234][12] = 8'd30;
        rom[234][13] = -8'd40;
        rom[234][14] = -8'd13;
        rom[234][15] = -8'd17;
        rom[234][16] = 8'd14;
        rom[234][17] = 8'd9;
        rom[234][18] = 8'd41;
        rom[234][19] = -8'd15;
        rom[234][20] = -8'd13;
        rom[234][21] = 8'd30;
        rom[234][22] = 8'd29;
        rom[234][23] = 8'd26;
        rom[234][24] = 8'd26;
        rom[234][25] = -8'd55;
        rom[234][26] = -8'd11;
        rom[234][27] = -8'd71;
        rom[234][28] = -8'd20;
        rom[234][29] = 8'd4;
        rom[234][30] = -8'd17;
        rom[234][31] = 8'd1;
        rom[235][0] = 8'd0;
        rom[235][1] = 8'd15;
        rom[235][2] = 8'd7;
        rom[235][3] = 8'd16;
        rom[235][4] = 8'd5;
        rom[235][5] = 8'd19;
        rom[235][6] = 8'd21;
        rom[235][7] = 8'd15;
        rom[235][8] = -8'd4;
        rom[235][9] = 8'd16;
        rom[235][10] = 8'd0;
        rom[235][11] = 8'd18;
        rom[235][12] = -8'd7;
        rom[235][13] = 8'd6;
        rom[235][14] = 8'd2;
        rom[235][15] = 8'd18;
        rom[235][16] = -8'd26;
        rom[235][17] = -8'd14;
        rom[235][18] = -8'd14;
        rom[235][19] = -8'd11;
        rom[235][20] = 8'd4;
        rom[235][21] = 8'd14;
        rom[235][22] = 8'd8;
        rom[235][23] = 8'd25;
        rom[235][24] = 8'd41;
        rom[235][25] = 8'd19;
        rom[235][26] = -8'd2;
        rom[235][27] = -8'd12;
        rom[235][28] = 8'd19;
        rom[235][29] = -8'd4;
        rom[235][30] = -8'd23;
        rom[235][31] = -8'd39;
        rom[236][0] = -8'd22;
        rom[236][1] = -8'd45;
        rom[236][2] = -8'd4;
        rom[236][3] = -8'd4;
        rom[236][4] = -8'd30;
        rom[236][5] = 8'd4;
        rom[236][6] = 8'd20;
        rom[236][7] = -8'd29;
        rom[236][8] = -8'd24;
        rom[236][9] = 8'd5;
        rom[236][10] = 8'd18;
        rom[236][11] = -8'd16;
        rom[236][12] = 8'd19;
        rom[236][13] = -8'd18;
        rom[236][14] = 8'd6;
        rom[236][15] = -8'd19;
        rom[236][16] = 8'd5;
        rom[236][17] = 8'd4;
        rom[236][18] = 8'd9;
        rom[236][19] = 8'd25;
        rom[236][20] = -8'd36;
        rom[236][21] = -8'd4;
        rom[236][22] = 8'd1;
        rom[236][23] = 8'd47;
        rom[236][24] = 8'd5;
        rom[236][25] = -8'd33;
        rom[236][26] = -8'd9;
        rom[236][27] = -8'd13;
        rom[236][28] = -8'd31;
        rom[236][29] = -8'd14;
        rom[236][30] = 8'd44;
        rom[236][31] = -8'd21;
        rom[237][0] = -8'd30;
        rom[237][1] = -8'd95;
        rom[237][2] = 8'd3;
        rom[237][3] = -8'd19;
        rom[237][4] = -8'd41;
        rom[237][5] = 8'd33;
        rom[237][6] = -8'd6;
        rom[237][7] = 8'd18;
        rom[237][8] = -8'd27;
        rom[237][9] = -8'd17;
        rom[237][10] = -8'd5;
        rom[237][11] = -8'd22;
        rom[237][12] = -8'd20;
        rom[237][13] = -8'd32;
        rom[237][14] = -8'd21;
        rom[237][15] = -8'd33;
        rom[237][16] = -8'd21;
        rom[237][17] = -8'd43;
        rom[237][18] = -8'd38;
        rom[237][19] = 8'd19;
        rom[237][20] = 8'd2;
        rom[237][21] = -8'd18;
        rom[237][22] = -8'd6;
        rom[237][23] = -8'd5;
        rom[237][24] = 8'd40;
        rom[237][25] = -8'd36;
        rom[237][26] = 8'd2;
        rom[237][27] = -8'd25;
        rom[237][28] = 8'd4;
        rom[237][29] = 8'd5;
        rom[237][30] = 8'd22;
        rom[237][31] = 8'd12;
        rom[238][0] = 8'd23;
        rom[238][1] = 8'd8;
        rom[238][2] = -8'd20;
        rom[238][3] = -8'd27;
        rom[238][4] = -8'd12;
        rom[238][5] = 8'd5;
        rom[238][6] = -8'd71;
        rom[238][7] = 8'd6;
        rom[238][8] = -8'd8;
        rom[238][9] = -8'd18;
        rom[238][10] = -8'd26;
        rom[238][11] = -8'd40;
        rom[238][12] = -8'd31;
        rom[238][13] = 8'd5;
        rom[238][14] = -8'd22;
        rom[238][15] = -8'd11;
        rom[238][16] = -8'd28;
        rom[238][17] = -8'd6;
        rom[238][18] = -8'd4;
        rom[238][19] = 8'd1;
        rom[238][20] = 8'd23;
        rom[238][21] = 8'd3;
        rom[238][22] = 8'd3;
        rom[238][23] = -8'd49;
        rom[238][24] = -8'd38;
        rom[238][25] = -8'd7;
        rom[238][26] = 8'd12;
        rom[238][27] = 8'd10;
        rom[238][28] = -8'd9;
        rom[238][29] = -8'd12;
        rom[238][30] = 8'd15;
        rom[238][31] = 8'd13;
        rom[239][0] = -8'd36;
        rom[239][1] = 8'd7;
        rom[239][2] = -8'd29;
        rom[239][3] = -8'd23;
        rom[239][4] = 8'd8;
        rom[239][5] = 8'd19;
        rom[239][6] = -8'd5;
        rom[239][7] = -8'd24;
        rom[239][8] = 8'd21;
        rom[239][9] = -8'd45;
        rom[239][10] = -8'd12;
        rom[239][11] = 8'd20;
        rom[239][12] = -8'd12;
        rom[239][13] = 8'd3;
        rom[239][14] = 8'd8;
        rom[239][15] = -8'd49;
        rom[239][16] = 8'd16;
        rom[239][17] = -8'd13;
        rom[239][18] = -8'd11;
        rom[239][19] = -8'd15;
        rom[239][20] = -8'd39;
        rom[239][21] = -8'd58;
        rom[239][22] = -8'd20;
        rom[239][23] = -8'd4;
        rom[239][24] = -8'd31;
        rom[239][25] = -8'd18;
        rom[239][26] = -8'd15;
        rom[239][27] = -8'd11;
        rom[239][28] = -8'd20;
        rom[239][29] = -8'd4;
        rom[239][30] = 8'd1;
        rom[239][31] = 8'd9;
        rom[240][0] = -8'd7;
        rom[240][1] = -8'd23;
        rom[240][2] = -8'd8;
        rom[240][3] = -8'd11;
        rom[240][4] = -8'd19;
        rom[240][5] = 8'd4;
        rom[240][6] = -8'd8;
        rom[240][7] = -8'd9;
        rom[240][8] = 8'd2;
        rom[240][9] = -8'd32;
        rom[240][10] = 8'd48;
        rom[240][11] = -8'd2;
        rom[240][12] = -8'd20;
        rom[240][13] = -8'd22;
        rom[240][14] = 8'd20;
        rom[240][15] = -8'd45;
        rom[240][16] = -8'd14;
        rom[240][17] = 8'd34;
        rom[240][18] = 8'd18;
        rom[240][19] = -8'd97;
        rom[240][20] = -8'd48;
        rom[240][21] = -8'd49;
        rom[240][22] = 8'd17;
        rom[240][23] = 8'd8;
        rom[240][24] = -8'd16;
        rom[240][25] = -8'd62;
        rom[240][26] = -8'd21;
        rom[240][27] = -8'd28;
        rom[240][28] = -8'd37;
        rom[240][29] = -8'd10;
        rom[240][30] = -8'd53;
        rom[240][31] = -8'd22;
        rom[241][0] = -8'd7;
        rom[241][1] = -8'd10;
        rom[241][2] = -8'd18;
        rom[241][3] = -8'd39;
        rom[241][4] = -8'd22;
        rom[241][5] = 8'd7;
        rom[241][6] = -8'd30;
        rom[241][7] = -8'd32;
        rom[241][8] = -8'd8;
        rom[241][9] = -8'd14;
        rom[241][10] = -8'd9;
        rom[241][11] = -8'd6;
        rom[241][12] = -8'd6;
        rom[241][13] = 8'd12;
        rom[241][14] = -8'd22;
        rom[241][15] = 8'd11;
        rom[241][16] = 8'd30;
        rom[241][17] = -8'd8;
        rom[241][18] = -8'd36;
        rom[241][19] = 8'd1;
        rom[241][20] = 8'd22;
        rom[241][21] = -8'd24;
        rom[241][22] = -8'd8;
        rom[241][23] = -8'd14;
        rom[241][24] = -8'd4;
        rom[241][25] = 8'd4;
        rom[241][26] = 8'd2;
        rom[241][27] = 8'd0;
        rom[241][28] = 8'd6;
        rom[241][29] = -8'd9;
        rom[241][30] = -8'd17;
        rom[241][31] = 8'd6;
        rom[242][0] = -8'd16;
        rom[242][1] = -8'd47;
        rom[242][2] = 8'd18;
        rom[242][3] = 8'd3;
        rom[242][4] = -8'd27;
        rom[242][5] = 8'd2;
        rom[242][6] = -8'd22;
        rom[242][7] = 8'd16;
        rom[242][8] = 8'd4;
        rom[242][9] = -8'd20;
        rom[242][10] = -8'd26;
        rom[242][11] = 8'd4;
        rom[242][12] = 8'd5;
        rom[242][13] = -8'd38;
        rom[242][14] = 8'd35;
        rom[242][15] = -8'd2;
        rom[242][16] = -8'd27;
        rom[242][17] = 8'd10;
        rom[242][18] = 8'd15;
        rom[242][19] = 8'd17;
        rom[242][20] = 8'd19;
        rom[242][21] = -8'd27;
        rom[242][22] = -8'd34;
        rom[242][23] = -8'd23;
        rom[242][24] = -8'd67;
        rom[242][25] = -8'd19;
        rom[242][26] = 8'd7;
        rom[242][27] = -8'd10;
        rom[242][28] = 8'd2;
        rom[242][29] = -8'd4;
        rom[242][30] = -8'd4;
        rom[242][31] = 8'd27;
        rom[243][0] = -8'd27;
        rom[243][1] = -8'd18;
        rom[243][2] = -8'd18;
        rom[243][3] = 8'd17;
        rom[243][4] = -8'd22;
        rom[243][5] = 8'd12;
        rom[243][6] = -8'd12;
        rom[243][7] = -8'd39;
        rom[243][8] = -8'd33;
        rom[243][9] = 8'd18;
        rom[243][10] = -8'd31;
        rom[243][11] = -8'd29;
        rom[243][12] = 8'd11;
        rom[243][13] = -8'd28;
        rom[243][14] = -8'd11;
        rom[243][15] = 8'd11;
        rom[243][16] = -8'd39;
        rom[243][17] = 8'd12;
        rom[243][18] = 8'd12;
        rom[243][19] = -8'd1;
        rom[243][20] = 8'd9;
        rom[243][21] = 8'd17;
        rom[243][22] = 8'd3;
        rom[243][23] = -8'd41;
        rom[243][24] = 8'd12;
        rom[243][25] = -8'd28;
        rom[243][26] = 8'd1;
        rom[243][27] = -8'd21;
        rom[243][28] = -8'd26;
        rom[243][29] = -8'd9;
        rom[243][30] = 8'd24;
        rom[243][31] = -8'd38;
        rom[244][0] = 8'd13;
        rom[244][1] = 8'd21;
        rom[244][2] = -8'd38;
        rom[244][3] = -8'd4;
        rom[244][4] = 8'd32;
        rom[244][5] = 8'd4;
        rom[244][6] = -8'd7;
        rom[244][7] = -8'd6;
        rom[244][8] = 8'd26;
        rom[244][9] = -8'd14;
        rom[244][10] = 8'd0;
        rom[244][11] = 8'd38;
        rom[244][12] = -8'd2;
        rom[244][13] = 8'd28;
        rom[244][14] = -8'd56;
        rom[244][15] = -8'd10;
        rom[244][16] = 8'd6;
        rom[244][17] = 8'd3;
        rom[244][18] = 8'd11;
        rom[244][19] = -8'd46;
        rom[244][20] = 8'd6;
        rom[244][21] = 8'd26;
        rom[244][22] = 8'd7;
        rom[244][23] = 8'd20;
        rom[244][24] = 8'd36;
        rom[244][25] = 8'd0;
        rom[244][26] = -8'd16;
        rom[244][27] = -8'd15;
        rom[244][28] = -8'd40;
        rom[244][29] = -8'd2;
        rom[244][30] = -8'd40;
        rom[244][31] = -8'd41;
        rom[245][0] = -8'd1;
        rom[245][1] = -8'd13;
        rom[245][2] = -8'd56;
        rom[245][3] = -8'd21;
        rom[245][4] = 8'd53;
        rom[245][5] = 8'd10;
        rom[245][6] = -8'd17;
        rom[245][7] = 8'd10;
        rom[245][8] = -8'd23;
        rom[245][9] = 8'd27;
        rom[245][10] = -8'd6;
        rom[245][11] = -8'd34;
        rom[245][12] = 8'd1;
        rom[245][13] = 8'd20;
        rom[245][14] = 8'd12;
        rom[245][15] = -8'd12;
        rom[245][16] = -8'd1;
        rom[245][17] = 8'd5;
        rom[245][18] = -8'd31;
        rom[245][19] = 8'd5;
        rom[245][20] = -8'd6;
        rom[245][21] = 8'd10;
        rom[245][22] = 8'd16;
        rom[245][23] = 8'd33;
        rom[245][24] = 8'd56;
        rom[245][25] = -8'd2;
        rom[245][26] = -8'd6;
        rom[245][27] = 8'd15;
        rom[245][28] = 8'd25;
        rom[245][29] = 8'd4;
        rom[245][30] = -8'd22;
        rom[245][31] = -8'd34;
        rom[246][0] = -8'd19;
        rom[246][1] = -8'd44;
        rom[246][2] = -8'd20;
        rom[246][3] = 8'd6;
        rom[246][4] = -8'd6;
        rom[246][5] = -8'd7;
        rom[246][6] = 8'd13;
        rom[246][7] = 8'd24;
        rom[246][8] = -8'd2;
        rom[246][9] = -8'd1;
        rom[246][10] = 8'd12;
        rom[246][11] = -8'd17;
        rom[246][12] = -8'd17;
        rom[246][13] = 8'd14;
        rom[246][14] = -8'd4;
        rom[246][15] = -8'd7;
        rom[246][16] = -8'd2;
        rom[246][17] = -8'd46;
        rom[246][18] = 8'd8;
        rom[246][19] = -8'd1;
        rom[246][20] = 8'd12;
        rom[246][21] = -8'd3;
        rom[246][22] = 8'd30;
        rom[246][23] = -8'd35;
        rom[246][24] = -8'd31;
        rom[246][25] = -8'd44;
        rom[246][26] = -8'd25;
        rom[246][27] = 8'd1;
        rom[246][28] = 8'd16;
        rom[246][29] = -8'd8;
        rom[246][30] = 8'd6;
        rom[246][31] = -8'd27;
        rom[247][0] = 8'd21;
        rom[247][1] = 8'd9;
        rom[247][2] = -8'd42;
        rom[247][3] = 8'd1;
        rom[247][4] = 8'd0;
        rom[247][5] = 8'd41;
        rom[247][6] = -8'd39;
        rom[247][7] = -8'd24;
        rom[247][8] = -8'd8;
        rom[247][9] = 8'd5;
        rom[247][10] = -8'd33;
        rom[247][11] = -8'd7;
        rom[247][12] = 8'd30;
        rom[247][13] = -8'd24;
        rom[247][14] = -8'd16;
        rom[247][15] = -8'd12;
        rom[247][16] = -8'd10;
        rom[247][17] = -8'd28;
        rom[247][18] = -8'd17;
        rom[247][19] = -8'd23;
        rom[247][20] = -8'd1;
        rom[247][21] = 8'd15;
        rom[247][22] = -8'd61;
        rom[247][23] = -8'd1;
        rom[247][24] = -8'd3;
        rom[247][25] = 8'd43;
        rom[247][26] = -8'd2;
        rom[247][27] = -8'd6;
        rom[247][28] = -8'd12;
        rom[247][29] = -8'd1;
        rom[247][30] = -8'd11;
        rom[247][31] = 8'd46;
        rom[248][0] = 8'd11;
        rom[248][1] = -8'd15;
        rom[248][2] = 8'd38;
        rom[248][3] = 8'd40;
        rom[248][4] = -8'd2;
        rom[248][5] = 8'd42;
        rom[248][6] = 8'd5;
        rom[248][7] = -8'd1;
        rom[248][8] = -8'd10;
        rom[248][9] = -8'd14;
        rom[248][10] = -8'd29;
        rom[248][11] = -8'd52;
        rom[248][12] = -8'd29;
        rom[248][13] = 8'd12;
        rom[248][14] = 8'd63;
        rom[248][15] = 8'd2;
        rom[248][16] = -8'd17;
        rom[248][17] = -8'd27;
        rom[248][18] = 8'd20;
        rom[248][19] = -8'd17;
        rom[248][20] = 8'd45;
        rom[248][21] = 8'd31;
        rom[248][22] = -8'd84;
        rom[248][23] = 8'd23;
        rom[248][24] = 8'd27;
        rom[248][25] = -8'd16;
        rom[248][26] = -8'd47;
        rom[248][27] = 8'd14;
        rom[248][28] = -8'd18;
        rom[248][29] = -8'd14;
        rom[248][30] = -8'd51;
        rom[248][31] = -8'd41;
        rom[249][0] = -8'd7;
        rom[249][1] = 8'd26;
        rom[249][2] = -8'd12;
        rom[249][3] = -8'd8;
        rom[249][4] = 8'd1;
        rom[249][5] = 8'd15;
        rom[249][6] = -8'd26;
        rom[249][7] = 8'd2;
        rom[249][8] = 8'd8;
        rom[249][9] = 8'd17;
        rom[249][10] = 8'd20;
        rom[249][11] = -8'd41;
        rom[249][12] = -8'd3;
        rom[249][13] = 8'd18;
        rom[249][14] = 8'd29;
        rom[249][15] = 8'd24;
        rom[249][16] = 8'd3;
        rom[249][17] = 8'd23;
        rom[249][18] = -8'd6;
        rom[249][19] = -8'd15;
        rom[249][20] = 8'd0;
        rom[249][21] = 8'd20;
        rom[249][22] = 8'd14;
        rom[249][23] = -8'd3;
        rom[249][24] = 8'd18;
        rom[249][25] = -8'd22;
        rom[249][26] = -8'd13;
        rom[249][27] = 8'd14;
        rom[249][28] = 8'd6;
        rom[249][29] = 8'd5;
        rom[249][30] = -8'd35;
        rom[249][31] = -8'd4;
        rom[250][0] = -8'd50;
        rom[250][1] = -8'd7;
        rom[250][2] = 8'd23;
        rom[250][3] = -8'd16;
        rom[250][4] = 8'd17;
        rom[250][5] = 8'd23;
        rom[250][6] = 8'd11;
        rom[250][7] = 8'd16;
        rom[250][8] = 8'd2;
        rom[250][9] = 8'd15;
        rom[250][10] = -8'd2;
        rom[250][11] = -8'd28;
        rom[250][12] = 8'd3;
        rom[250][13] = -8'd6;
        rom[250][14] = -8'd6;
        rom[250][15] = 8'd12;
        rom[250][16] = 8'd30;
        rom[250][17] = -8'd23;
        rom[250][18] = 8'd12;
        rom[250][19] = 8'd16;
        rom[250][20] = 8'd5;
        rom[250][21] = -8'd18;
        rom[250][22] = -8'd20;
        rom[250][23] = 8'd7;
        rom[250][24] = -8'd32;
        rom[250][25] = 8'd17;
        rom[250][26] = 8'd3;
        rom[250][27] = -8'd32;
        rom[250][28] = -8'd10;
        rom[250][29] = -8'd4;
        rom[250][30] = -8'd2;
        rom[250][31] = -8'd7;
        rom[251][0] = 8'd23;
        rom[251][1] = 8'd19;
        rom[251][2] = -8'd8;
        rom[251][3] = 8'd2;
        rom[251][4] = -8'd15;
        rom[251][5] = -8'd8;
        rom[251][6] = -8'd5;
        rom[251][7] = -8'd9;
        rom[251][8] = -8'd2;
        rom[251][9] = -8'd2;
        rom[251][10] = -8'd12;
        rom[251][11] = 8'd34;
        rom[251][12] = -8'd52;
        rom[251][13] = 8'd4;
        rom[251][14] = 8'd6;
        rom[251][15] = -8'd11;
        rom[251][16] = 8'd9;
        rom[251][17] = -8'd4;
        rom[251][18] = -8'd11;
        rom[251][19] = 8'd11;
        rom[251][20] = 8'd48;
        rom[251][21] = 8'd16;
        rom[251][22] = -8'd18;
        rom[251][23] = -8'd9;
        rom[251][24] = -8'd16;
        rom[251][25] = 8'd2;
        rom[251][26] = -8'd2;
        rom[251][27] = 8'd10;
        rom[251][28] = 8'd7;
        rom[251][29] = -8'd5;
        rom[251][30] = 8'd7;
        rom[251][31] = 8'd7;
        rom[252][0] = -8'd31;
        rom[252][1] = -8'd9;
        rom[252][2] = 8'd6;
        rom[252][3] = 8'd0;
        rom[252][4] = -8'd15;
        rom[252][5] = -8'd19;
        rom[252][6] = -8'd1;
        rom[252][7] = 8'd15;
        rom[252][8] = 8'd2;
        rom[252][9] = 8'd5;
        rom[252][10] = -8'd17;
        rom[252][11] = 8'd14;
        rom[252][12] = -8'd23;
        rom[252][13] = -8'd37;
        rom[252][14] = 8'd17;
        rom[252][15] = -8'd27;
        rom[252][16] = -8'd10;
        rom[252][17] = -8'd12;
        rom[252][18] = 8'd32;
        rom[252][19] = -8'd24;
        rom[252][20] = -8'd51;
        rom[252][21] = 8'd19;
        rom[252][22] = 8'd13;
        rom[252][23] = 8'd41;
        rom[252][24] = 8'd14;
        rom[252][25] = 8'd5;
        rom[252][26] = -8'd1;
        rom[252][27] = -8'd58;
        rom[252][28] = 8'd12;
        rom[252][29] = 8'd1;
        rom[252][30] = -8'd3;
        rom[252][31] = -8'd45;
        rom[253][0] = 8'd7;
        rom[253][1] = 8'd23;
        rom[253][2] = -8'd19;
        rom[253][3] = -8'd5;
        rom[253][4] = -8'd35;
        rom[253][5] = -8'd5;
        rom[253][6] = 8'd35;
        rom[253][7] = -8'd45;
        rom[253][8] = -8'd7;
        rom[253][9] = -8'd16;
        rom[253][10] = -8'd24;
        rom[253][11] = -8'd47;
        rom[253][12] = -8'd64;
        rom[253][13] = 8'd1;
        rom[253][14] = 8'd4;
        rom[253][15] = -8'd3;
        rom[253][16] = 8'd10;
        rom[253][17] = 8'd25;
        rom[253][18] = 8'd20;
        rom[253][19] = -8'd15;
        rom[253][20] = 8'd47;
        rom[253][21] = 8'd8;
        rom[253][22] = 8'd13;
        rom[253][23] = 8'd9;
        rom[253][24] = 8'd25;
        rom[253][25] = -8'd17;
        rom[253][26] = -8'd24;
        rom[253][27] = -8'd13;
        rom[253][28] = 8'd4;
        rom[253][29] = -8'd11;
        rom[253][30] = 8'd26;
        rom[253][31] = -8'd13;
        rom[254][0] = -8'd5;
        rom[254][1] = 8'd9;
        rom[254][2] = 8'd19;
        rom[254][3] = -8'd36;
        rom[254][4] = 8'd1;
        rom[254][5] = 8'd2;
        rom[254][6] = -8'd9;
        rom[254][7] = -8'd25;
        rom[254][8] = -8'd4;
        rom[254][9] = -8'd7;
        rom[254][10] = 8'd0;
        rom[254][11] = 8'd37;
        rom[254][12] = -8'd42;
        rom[254][13] = -8'd4;
        rom[254][14] = 8'd9;
        rom[254][15] = 8'd24;
        rom[254][16] = 8'd34;
        rom[254][17] = 8'd8;
        rom[254][18] = 8'd40;
        rom[254][19] = -8'd18;
        rom[254][20] = -8'd2;
        rom[254][21] = 8'd7;
        rom[254][22] = 8'd50;
        rom[254][23] = 8'd34;
        rom[254][24] = 8'd42;
        rom[254][25] = 8'd14;
        rom[254][26] = -8'd2;
        rom[254][27] = 8'd17;
        rom[254][28] = 8'd11;
        rom[254][29] = 8'd9;
        rom[254][30] = -8'd6;
        rom[254][31] = -8'd36;
        rom[255][0] = 8'd2;
        rom[255][1] = -8'd1;
        rom[255][2] = 8'd60;
        rom[255][3] = -8'd6;
        rom[255][4] = -8'd9;
        rom[255][5] = -8'd14;
        rom[255][6] = -8'd61;
        rom[255][7] = 8'd13;
        rom[255][8] = 8'd7;
        rom[255][9] = -8'd22;
        rom[255][10] = -8'd5;
        rom[255][11] = -8'd7;
        rom[255][12] = 8'd36;
        rom[255][13] = -8'd55;
        rom[255][14] = -8'd12;
        rom[255][15] = -8'd17;
        rom[255][16] = -8'd25;
        rom[255][17] = -8'd34;
        rom[255][18] = 8'd7;
        rom[255][19] = -8'd7;
        rom[255][20] = -8'd43;
        rom[255][21] = 8'd0;
        rom[255][22] = -8'd36;
        rom[255][23] = -8'd41;
        rom[255][24] = 8'd9;
        rom[255][25] = 8'd25;
        rom[255][26] = -8'd19;
        rom[255][27] = 8'd12;
        rom[255][28] = -8'd6;
        rom[255][29] = 8'd9;
        rom[255][30] = -8'd31;
        rom[255][31] = -8'd32;
        rom[256][0] = 8'd11;
        rom[256][1] = -8'd49;
        rom[256][2] = -8'd33;
        rom[256][3] = -8'd13;
        rom[256][4] = -8'd4;
        rom[256][5] = 8'd9;
        rom[256][6] = -8'd31;
        rom[256][7] = -8'd23;
        rom[256][8] = -8'd11;
        rom[256][9] = 8'd21;
        rom[256][10] = 8'd29;
        rom[256][11] = 8'd6;
        rom[256][12] = -8'd45;
        rom[256][13] = 8'd21;
        rom[256][14] = 8'd14;
        rom[256][15] = -8'd24;
        rom[256][16] = -8'd5;
        rom[256][17] = 8'd11;
        rom[256][18] = -8'd13;
        rom[256][19] = -8'd18;
        rom[256][20] = 8'd12;
        rom[256][21] = -8'd12;
        rom[256][22] = 8'd26;
        rom[256][23] = 8'd4;
        rom[256][24] = -8'd5;
        rom[256][25] = 8'd5;
        rom[256][26] = -8'd9;
        rom[256][27] = 8'd20;
        rom[256][28] = 8'd10;
        rom[256][29] = -8'd9;
        rom[256][30] = 8'd27;
        rom[256][31] = -8'd13;
        rom[257][0] = -8'd13;
        rom[257][1] = 8'd24;
        rom[257][2] = 8'd26;
        rom[257][3] = 8'd31;
        rom[257][4] = -8'd42;
        rom[257][5] = -8'd6;
        rom[257][6] = 8'd15;
        rom[257][7] = 8'd52;
        rom[257][8] = 8'd31;
        rom[257][9] = 8'd37;
        rom[257][10] = -8'd11;
        rom[257][11] = 8'd21;
        rom[257][12] = 8'd26;
        rom[257][13] = -8'd35;
        rom[257][14] = 8'd3;
        rom[257][15] = -8'd21;
        rom[257][16] = -8'd8;
        rom[257][17] = 8'd5;
        rom[257][18] = 8'd23;
        rom[257][19] = -8'd9;
        rom[257][20] = 8'd13;
        rom[257][21] = -8'd2;
        rom[257][22] = 8'd50;
        rom[257][23] = 8'd3;
        rom[257][24] = 8'd6;
        rom[257][25] = 8'd34;
        rom[257][26] = 8'd6;
        rom[257][27] = -8'd50;
        rom[257][28] = -8'd1;
        rom[257][29] = -8'd17;
        rom[257][30] = -8'd39;
        rom[257][31] = 8'd38;
        rom[258][0] = 8'd12;
        rom[258][1] = 8'd17;
        rom[258][2] = -8'd44;
        rom[258][3] = 8'd38;
        rom[258][4] = -8'd12;
        rom[258][5] = 8'd24;
        rom[258][6] = 8'd40;
        rom[258][7] = -8'd11;
        rom[258][8] = -8'd38;
        rom[258][9] = -8'd31;
        rom[258][10] = -8'd46;
        rom[258][11] = -8'd6;
        rom[258][12] = 8'd23;
        rom[258][13] = -8'd50;
        rom[258][14] = -8'd34;
        rom[258][15] = -8'd18;
        rom[258][16] = 8'd12;
        rom[258][17] = 8'd6;
        rom[258][18] = -8'd28;
        rom[258][19] = -8'd12;
        rom[258][20] = -8'd64;
        rom[258][21] = 8'd34;
        rom[258][22] = -8'd30;
        rom[258][23] = 8'd47;
        rom[258][24] = -8'd33;
        rom[258][25] = -8'd10;
        rom[258][26] = 8'd28;
        rom[258][27] = 8'd38;
        rom[258][28] = 8'd41;
        rom[258][29] = -8'd6;
        rom[258][30] = -8'd15;
        rom[258][31] = 8'd6;
        rom[259][0] = 8'd25;
        rom[259][1] = -8'd47;
        rom[259][2] = -8'd17;
        rom[259][3] = 8'd5;
        rom[259][4] = -8'd66;
        rom[259][5] = -8'd18;
        rom[259][6] = -8'd23;
        rom[259][7] = -8'd8;
        rom[259][8] = 8'd19;
        rom[259][9] = 8'd4;
        rom[259][10] = -8'd46;
        rom[259][11] = 8'd21;
        rom[259][12] = -8'd71;
        rom[259][13] = 8'd25;
        rom[259][14] = -8'd31;
        rom[259][15] = -8'd9;
        rom[259][16] = 8'd18;
        rom[259][17] = 8'd13;
        rom[259][18] = -8'd3;
        rom[259][19] = -8'd23;
        rom[259][20] = 8'd6;
        rom[259][21] = -8'd35;
        rom[259][22] = 8'd11;
        rom[259][23] = 8'd9;
        rom[259][24] = -8'd16;
        rom[259][25] = -8'd23;
        rom[259][26] = 8'd37;
        rom[259][27] = 8'd27;
        rom[259][28] = -8'd60;
        rom[259][29] = 8'd11;
        rom[259][30] = 8'd33;
        rom[259][31] = -8'd17;
        rom[260][0] = 8'd4;
        rom[260][1] = -8'd6;
        rom[260][2] = 8'd8;
        rom[260][3] = -8'd4;
        rom[260][4] = -8'd48;
        rom[260][5] = -8'd26;
        rom[260][6] = 8'd9;
        rom[260][7] = 8'd30;
        rom[260][8] = 8'd2;
        rom[260][9] = 8'd22;
        rom[260][10] = 8'd4;
        rom[260][11] = -8'd24;
        rom[260][12] = 8'd8;
        rom[260][13] = 8'd6;
        rom[260][14] = 8'd44;
        rom[260][15] = 8'd36;
        rom[260][16] = 8'd4;
        rom[260][17] = 8'd24;
        rom[260][18] = 8'd11;
        rom[260][19] = 8'd1;
        rom[260][20] = 8'd2;
        rom[260][21] = -8'd11;
        rom[260][22] = -8'd6;
        rom[260][23] = -8'd7;
        rom[260][24] = 8'd34;
        rom[260][25] = -8'd26;
        rom[260][26] = -8'd16;
        rom[260][27] = -8'd29;
        rom[260][28] = 8'd7;
        rom[260][29] = 8'd9;
        rom[260][30] = 8'd27;
        rom[260][31] = -8'd11;
        rom[261][0] = 8'd1;
        rom[261][1] = -8'd5;
        rom[261][2] = -8'd25;
        rom[261][3] = -8'd17;
        rom[261][4] = 8'd77;
        rom[261][5] = -8'd3;
        rom[261][6] = 8'd48;
        rom[261][7] = -8'd18;
        rom[261][8] = 8'd12;
        rom[261][9] = -8'd6;
        rom[261][10] = -8'd29;
        rom[261][11] = -8'd19;
        rom[261][12] = 8'd19;
        rom[261][13] = 8'd28;
        rom[261][14] = 8'd6;
        rom[261][15] = -8'd21;
        rom[261][16] = 8'd41;
        rom[261][17] = 8'd10;
        rom[261][18] = -8'd30;
        rom[261][19] = -8'd3;
        rom[261][20] = -8'd31;
        rom[261][21] = 8'd37;
        rom[261][22] = 8'd13;
        rom[261][23] = 8'd6;
        rom[261][24] = -8'd14;
        rom[261][25] = -8'd53;
        rom[261][26] = -8'd23;
        rom[261][27] = 8'd0;
        rom[261][28] = 8'd26;
        rom[261][29] = -8'd9;
        rom[261][30] = -8'd61;
        rom[261][31] = 8'd3;
        rom[262][0] = -8'd24;
        rom[262][1] = 8'd21;
        rom[262][2] = 8'd35;
        rom[262][3] = -8'd16;
        rom[262][4] = -8'd7;
        rom[262][5] = 8'd8;
        rom[262][6] = -8'd66;
        rom[262][7] = -8'd15;
        rom[262][8] = -8'd31;
        rom[262][9] = -8'd17;
        rom[262][10] = -8'd36;
        rom[262][11] = -8'd55;
        rom[262][12] = 8'd1;
        rom[262][13] = 8'd26;
        rom[262][14] = -8'd6;
        rom[262][15] = -8'd16;
        rom[262][16] = 8'd11;
        rom[262][17] = 8'd13;
        rom[262][18] = -8'd9;
        rom[262][19] = 8'd16;
        rom[262][20] = 8'd16;
        rom[262][21] = -8'd13;
        rom[262][22] = -8'd23;
        rom[262][23] = -8'd19;
        rom[262][24] = -8'd8;
        rom[262][25] = 8'd32;
        rom[262][26] = 8'd22;
        rom[262][27] = 8'd13;
        rom[262][28] = 8'd3;
        rom[262][29] = -8'd8;
        rom[262][30] = 8'd3;
        rom[262][31] = -8'd14;
        rom[263][0] = 8'd7;
        rom[263][1] = 8'd15;
        rom[263][2] = 8'd28;
        rom[263][3] = 8'd1;
        rom[263][4] = -8'd11;
        rom[263][5] = -8'd16;
        rom[263][6] = -8'd61;
        rom[263][7] = 8'd18;
        rom[263][8] = 8'd14;
        rom[263][9] = 8'd13;
        rom[263][10] = 8'd5;
        rom[263][11] = 8'd2;
        rom[263][12] = -8'd22;
        rom[263][13] = -8'd6;
        rom[263][14] = -8'd35;
        rom[263][15] = 8'd28;
        rom[263][16] = 8'd3;
        rom[263][17] = -8'd14;
        rom[263][18] = 8'd33;
        rom[263][19] = 8'd2;
        rom[263][20] = 8'd11;
        rom[263][21] = -8'd14;
        rom[263][22] = 8'd7;
        rom[263][23] = -8'd27;
        rom[263][24] = 8'd3;
        rom[263][25] = 8'd30;
        rom[263][26] = 8'd43;
        rom[263][27] = 8'd12;
        rom[263][28] = 8'd16;
        rom[263][29] = 8'd1;
        rom[263][30] = -8'd13;
        rom[263][31] = -8'd15;
        rom[264][0] = 8'd4;
        rom[264][1] = -8'd59;
        rom[264][2] = -8'd5;
        rom[264][3] = -8'd6;
        rom[264][4] = -8'd26;
        rom[264][5] = -8'd3;
        rom[264][6] = -8'd70;
        rom[264][7] = -8'd3;
        rom[264][8] = 8'd12;
        rom[264][9] = 8'd1;
        rom[264][10] = 8'd30;
        rom[264][11] = 8'd30;
        rom[264][12] = -8'd5;
        rom[264][13] = -8'd27;
        rom[264][14] = -8'd9;
        rom[264][15] = -8'd11;
        rom[264][16] = -8'd26;
        rom[264][17] = 8'd16;
        rom[264][18] = 8'd2;
        rom[264][19] = 8'd5;
        rom[264][20] = -8'd32;
        rom[264][21] = -8'd23;
        rom[264][22] = 8'd3;
        rom[264][23] = -8'd1;
        rom[264][24] = -8'd13;
        rom[264][25] = -8'd23;
        rom[264][26] = 8'd2;
        rom[264][27] = -8'd17;
        rom[264][28] = -8'd12;
        rom[264][29] = -8'd13;
        rom[264][30] = -8'd50;
        rom[264][31] = -8'd6;
        rom[265][0] = 8'd23;
        rom[265][1] = -8'd32;
        rom[265][2] = -8'd13;
        rom[265][3] = -8'd4;
        rom[265][4] = -8'd23;
        rom[265][5] = -8'd10;
        rom[265][6] = -8'd7;
        rom[265][7] = 8'd7;
        rom[265][8] = -8'd25;
        rom[265][9] = 8'd4;
        rom[265][10] = -8'd50;
        rom[265][11] = -8'd13;
        rom[265][12] = -8'd15;
        rom[265][13] = -8'd8;
        rom[265][14] = -8'd23;
        rom[265][15] = 8'd52;
        rom[265][16] = 8'd28;
        rom[265][17] = -8'd9;
        rom[265][18] = -8'd18;
        rom[265][19] = -8'd32;
        rom[265][20] = 8'd25;
        rom[265][21] = -8'd39;
        rom[265][22] = -8'd11;
        rom[265][23] = 8'd25;
        rom[265][24] = 8'd11;
        rom[265][25] = -8'd34;
        rom[265][26] = -8'd23;
        rom[265][27] = 8'd23;
        rom[265][28] = 8'd16;
        rom[265][29] = -8'd12;
        rom[265][30] = 8'd15;
        rom[265][31] = 8'd27;
        rom[266][0] = -8'd31;
        rom[266][1] = 8'd22;
        rom[266][2] = -8'd20;
        rom[266][3] = 8'd42;
        rom[266][4] = -8'd1;
        rom[266][5] = 8'd29;
        rom[266][6] = -8'd33;
        rom[266][7] = 8'd7;
        rom[266][8] = -8'd33;
        rom[266][9] = -8'd13;
        rom[266][10] = -8'd1;
        rom[266][11] = 8'd58;
        rom[266][12] = 8'd39;
        rom[266][13] = -8'd11;
        rom[266][14] = -8'd22;
        rom[266][15] = -8'd24;
        rom[266][16] = -8'd2;
        rom[266][17] = -8'd11;
        rom[266][18] = 8'd11;
        rom[266][19] = -8'd19;
        rom[266][20] = -8'd5;
        rom[266][21] = 8'd40;
        rom[266][22] = 8'd33;
        rom[266][23] = -8'd23;
        rom[266][24] = 8'd36;
        rom[266][25] = 8'd1;
        rom[266][26] = -8'd8;
        rom[266][27] = -8'd45;
        rom[266][28] = 8'd13;
        rom[266][29] = 8'd13;
        rom[266][30] = 8'd22;
        rom[266][31] = 8'd16;
        rom[267][0] = -8'd10;
        rom[267][1] = 8'd2;
        rom[267][2] = 8'd24;
        rom[267][3] = -8'd4;
        rom[267][4] = 8'd5;
        rom[267][5] = 8'd3;
        rom[267][6] = 8'd20;
        rom[267][7] = -8'd9;
        rom[267][8] = 8'd8;
        rom[267][9] = 8'd10;
        rom[267][10] = -8'd26;
        rom[267][11] = 8'd12;
        rom[267][12] = -8'd35;
        rom[267][13] = -8'd9;
        rom[267][14] = -8'd9;
        rom[267][15] = 8'd23;
        rom[267][16] = -8'd7;
        rom[267][17] = -8'd17;
        rom[267][18] = 8'd19;
        rom[267][19] = 8'd5;
        rom[267][20] = 8'd12;
        rom[267][21] = 8'd29;
        rom[267][22] = -8'd15;
        rom[267][23] = -8'd56;
        rom[267][24] = 8'd17;
        rom[267][25] = 8'd0;
        rom[267][26] = -8'd6;
        rom[267][27] = -8'd7;
        rom[267][28] = 8'd25;
        rom[267][29] = -8'd8;
        rom[267][30] = -8'd17;
        rom[267][31] = -8'd25;
        rom[268][0] = 8'd37;
        rom[268][1] = -8'd13;
        rom[268][2] = -8'd34;
        rom[268][3] = 8'd4;
        rom[268][4] = 8'd18;
        rom[268][5] = -8'd46;
        rom[268][6] = 8'd8;
        rom[268][7] = 8'd0;
        rom[268][8] = -8'd33;
        rom[268][9] = 8'd22;
        rom[268][10] = 8'd22;
        rom[268][11] = 8'd21;
        rom[268][12] = 8'd40;
        rom[268][13] = -8'd2;
        rom[268][14] = -8'd23;
        rom[268][15] = 8'd18;
        rom[268][16] = 8'd25;
        rom[268][17] = 8'd18;
        rom[268][18] = -8'd42;
        rom[268][19] = 8'd25;
        rom[268][20] = -8'd39;
        rom[268][21] = 8'd15;
        rom[268][22] = 8'd29;
        rom[268][23] = 8'd46;
        rom[268][24] = -8'd22;
        rom[268][25] = -8'd29;
        rom[268][26] = -8'd9;
        rom[268][27] = 8'd2;
        rom[268][28] = 8'd1;
        rom[268][29] = -8'd13;
        rom[268][30] = 8'd37;
        rom[268][31] = 8'd17;
        rom[269][0] = 8'd7;
        rom[269][1] = -8'd35;
        rom[269][2] = -8'd43;
        rom[269][3] = 8'd6;
        rom[269][4] = 8'd1;
        rom[269][5] = -8'd40;
        rom[269][6] = 8'd31;
        rom[269][7] = -8'd3;
        rom[269][8] = -8'd20;
        rom[269][9] = 8'd8;
        rom[269][10] = -8'd28;
        rom[269][11] = -8'd34;
        rom[269][12] = -8'd4;
        rom[269][13] = -8'd6;
        rom[269][14] = -8'd29;
        rom[269][15] = -8'd31;
        rom[269][16] = -8'd24;
        rom[269][17] = 8'd7;
        rom[269][18] = 8'd0;
        rom[269][19] = 8'd37;
        rom[269][20] = 8'd20;
        rom[269][21] = 8'd10;
        rom[269][22] = -8'd11;
        rom[269][23] = 8'd1;
        rom[269][24] = 8'd15;
        rom[269][25] = -8'd26;
        rom[269][26] = 8'd18;
        rom[269][27] = 8'd24;
        rom[269][28] = -8'd19;
        rom[269][29] = -8'd6;
        rom[269][30] = 8'd29;
        rom[269][31] = -8'd28;
        rom[270][0] = 8'd11;
        rom[270][1] = -8'd5;
        rom[270][2] = 8'd23;
        rom[270][3] = -8'd49;
        rom[270][4] = -8'd17;
        rom[270][5] = -8'd16;
        rom[270][6] = -8'd64;
        rom[270][7] = 8'd33;
        rom[270][8] = 8'd8;
        rom[270][9] = 8'd0;
        rom[270][10] = -8'd9;
        rom[270][11] = -8'd59;
        rom[270][12] = -8'd19;
        rom[270][13] = 8'd17;
        rom[270][14] = 8'd18;
        rom[270][15] = 8'd3;
        rom[270][16] = -8'd42;
        rom[270][17] = 8'd1;
        rom[270][18] = 8'd14;
        rom[270][19] = 8'd5;
        rom[270][20] = 8'd18;
        rom[270][21] = -8'd7;
        rom[270][22] = 8'd26;
        rom[270][23] = -8'd36;
        rom[270][24] = -8'd10;
        rom[270][25] = -8'd7;
        rom[270][26] = 8'd20;
        rom[270][27] = 8'd0;
        rom[270][28] = -8'd22;
        rom[270][29] = -8'd17;
        rom[270][30] = 8'd30;
        rom[270][31] = -8'd5;
        rom[271][0] = 8'd45;
        rom[271][1] = -8'd39;
        rom[271][2] = -8'd56;
        rom[271][3] = 8'd2;
        rom[271][4] = 8'd6;
        rom[271][5] = 8'd10;
        rom[271][6] = -8'd37;
        rom[271][7] = 8'd18;
        rom[271][8] = 8'd3;
        rom[271][9] = -8'd48;
        rom[271][10] = -8'd8;
        rom[271][11] = 8'd16;
        rom[271][12] = -8'd1;
        rom[271][13] = 8'd7;
        rom[271][14] = 8'd5;
        rom[271][15] = -8'd71;
        rom[271][16] = 8'd9;
        rom[271][17] = 8'd32;
        rom[271][18] = 8'd14;
        rom[271][19] = -8'd5;
        rom[271][20] = -8'd25;
        rom[271][21] = -8'd67;
        rom[271][22] = 8'd4;
        rom[271][23] = 8'd7;
        rom[271][24] = -8'd27;
        rom[271][25] = -8'd2;
        rom[271][26] = -8'd24;
        rom[271][27] = 8'd31;
        rom[271][28] = -8'd7;
        rom[271][29] = -8'd9;
        rom[271][30] = 8'd26;
        rom[271][31] = 8'd8;
        rom[272][0] = 8'd12;
        rom[272][1] = -8'd20;
        rom[272][2] = -8'd36;
        rom[272][3] = 8'd10;
        rom[272][4] = -8'd5;
        rom[272][5] = -8'd4;
        rom[272][6] = -8'd38;
        rom[272][7] = -8'd35;
        rom[272][8] = 8'd24;
        rom[272][9] = -8'd20;
        rom[272][10] = 8'd29;
        rom[272][11] = 8'd4;
        rom[272][12] = 8'd5;
        rom[272][13] = 8'd7;
        rom[272][14] = -8'd26;
        rom[272][15] = -8'd24;
        rom[272][16] = 8'd12;
        rom[272][17] = 8'd11;
        rom[272][18] = 8'd26;
        rom[272][19] = -8'd75;
        rom[272][20] = -8'd82;
        rom[272][21] = -8'd68;
        rom[272][22] = 8'd10;
        rom[272][23] = 8'd50;
        rom[272][24] = 8'd17;
        rom[272][25] = -8'd30;
        rom[272][26] = -8'd3;
        rom[272][27] = 8'd9;
        rom[272][28] = -8'd20;
        rom[272][29] = -8'd10;
        rom[272][30] = -8'd31;
        rom[272][31] = -8'd22;
        rom[273][0] = 8'd9;
        rom[273][1] = 8'd14;
        rom[273][2] = 8'd31;
        rom[273][3] = -8'd6;
        rom[273][4] = -8'd28;
        rom[273][5] = 8'd16;
        rom[273][6] = -8'd35;
        rom[273][7] = 8'd16;
        rom[273][8] = -8'd18;
        rom[273][9] = -8'd24;
        rom[273][10] = 8'd6;
        rom[273][11] = -8'd10;
        rom[273][12] = 8'd5;
        rom[273][13] = 8'd21;
        rom[273][14] = 8'd31;
        rom[273][15] = 8'd45;
        rom[273][16] = -8'd25;
        rom[273][17] = 8'd11;
        rom[273][18] = -8'd25;
        rom[273][19] = -8'd5;
        rom[273][20] = 8'd21;
        rom[273][21] = 8'd1;
        rom[273][22] = -8'd2;
        rom[273][23] = 8'd11;
        rom[273][24] = 8'd9;
        rom[273][25] = -8'd12;
        rom[273][26] = 8'd8;
        rom[273][27] = 8'd34;
        rom[273][28] = 8'd34;
        rom[273][29] = 8'd3;
        rom[273][30] = -8'd33;
        rom[273][31] = -8'd24;
        rom[274][0] = 8'd4;
        rom[274][1] = -8'd53;
        rom[274][2] = -8'd18;
        rom[274][3] = 8'd18;
        rom[274][4] = -8'd21;
        rom[274][5] = -8'd44;
        rom[274][6] = -8'd10;
        rom[274][7] = 8'd16;
        rom[274][8] = -8'd26;
        rom[274][9] = 8'd7;
        rom[274][10] = -8'd25;
        rom[274][11] = -8'd5;
        rom[274][12] = 8'd38;
        rom[274][13] = -8'd27;
        rom[274][14] = 8'd34;
        rom[274][15] = -8'd36;
        rom[274][16] = -8'd76;
        rom[274][17] = 8'd20;
        rom[274][18] = 8'd29;
        rom[274][19] = 8'd11;
        rom[274][20] = -8'd3;
        rom[274][21] = -8'd19;
        rom[274][22] = -8'd21;
        rom[274][23] = 8'd31;
        rom[274][24] = -8'd52;
        rom[274][25] = 8'd2;
        rom[274][26] = 8'd20;
        rom[274][27] = 8'd4;
        rom[274][28] = 8'd0;
        rom[274][29] = -8'd9;
        rom[274][30] = 8'd12;
        rom[274][31] = 8'd24;
        rom[275][0] = 8'd7;
        rom[275][1] = 8'd31;
        rom[275][2] = 8'd14;
        rom[275][3] = -8'd17;
        rom[275][4] = 8'd28;
        rom[275][5] = -8'd17;
        rom[275][6] = -8'd4;
        rom[275][7] = -8'd41;
        rom[275][8] = -8'd27;
        rom[275][9] = 8'd14;
        rom[275][10] = 8'd5;
        rom[275][11] = -8'd6;
        rom[275][12] = 8'd7;
        rom[275][13] = -8'd6;
        rom[275][14] = -8'd4;
        rom[275][15] = 8'd18;
        rom[275][16] = 8'd9;
        rom[275][17] = 8'd14;
        rom[275][18] = 8'd22;
        rom[275][19] = 8'd2;
        rom[275][20] = 8'd8;
        rom[275][21] = 8'd15;
        rom[275][22] = -8'd11;
        rom[275][23] = 8'd8;
        rom[275][24] = 8'd18;
        rom[275][25] = -8'd13;
        rom[275][26] = 8'd8;
        rom[275][27] = -8'd26;
        rom[275][28] = -8'd14;
        rom[275][29] = -8'd15;
        rom[275][30] = 8'd18;
        rom[275][31] = 8'd1;
        rom[276][0] = 8'd27;
        rom[276][1] = 8'd19;
        rom[276][2] = -8'd34;
        rom[276][3] = 8'd4;
        rom[276][4] = 8'd25;
        rom[276][5] = 8'd45;
        rom[276][6] = 8'd27;
        rom[276][7] = -8'd40;
        rom[276][8] = 8'd33;
        rom[276][9] = -8'd9;
        rom[276][10] = -8'd2;
        rom[276][11] = -8'd3;
        rom[276][12] = 8'd3;
        rom[276][13] = 8'd23;
        rom[276][14] = -8'd82;
        rom[276][15] = 8'd17;
        rom[276][16] = 8'd6;
        rom[276][17] = -8'd29;
        rom[276][18] = 8'd31;
        rom[276][19] = -8'd45;
        rom[276][20] = 8'd18;
        rom[276][21] = 8'd19;
        rom[276][22] = -8'd6;
        rom[276][23] = -8'd28;
        rom[276][24] = 8'd37;
        rom[276][25] = 8'd16;
        rom[276][26] = -8'd14;
        rom[276][27] = -8'd27;
        rom[276][28] = 8'd0;
        rom[276][29] = -8'd2;
        rom[276][30] = -8'd27;
        rom[276][31] = 8'd3;
        rom[277][0] = 8'd22;
        rom[277][1] = -8'd12;
        rom[277][2] = 8'd6;
        rom[277][3] = -8'd26;
        rom[277][4] = 8'd55;
        rom[277][5] = -8'd19;
        rom[277][6] = 8'd15;
        rom[277][7] = 8'd11;
        rom[277][8] = 8'd22;
        rom[277][9] = 8'd15;
        rom[277][10] = -8'd17;
        rom[277][11] = -8'd22;
        rom[277][12] = 8'd17;
        rom[277][13] = 8'd2;
        rom[277][14] = 8'd9;
        rom[277][15] = 8'd9;
        rom[277][16] = -8'd25;
        rom[277][17] = -8'd34;
        rom[277][18] = -8'd33;
        rom[277][19] = -8'd3;
        rom[277][20] = -8'd8;
        rom[277][21] = -8'd33;
        rom[277][22] = 8'd28;
        rom[277][23] = -8'd20;
        rom[277][24] = 8'd27;
        rom[277][25] = 8'd0;
        rom[277][26] = -8'd20;
        rom[277][27] = 8'd61;
        rom[277][28] = 8'd17;
        rom[277][29] = -8'd3;
        rom[277][30] = -8'd15;
        rom[277][31] = 8'd24;
        rom[278][0] = -8'd31;
        rom[278][1] = -8'd64;
        rom[278][2] = 8'd34;
        rom[278][3] = 8'd14;
        rom[278][4] = 8'd15;
        rom[278][5] = -8'd1;
        rom[278][6] = -8'd8;
        rom[278][7] = 8'd41;
        rom[278][8] = -8'd26;
        rom[278][9] = 8'd14;
        rom[278][10] = 8'd15;
        rom[278][11] = -8'd19;
        rom[278][12] = -8'd26;
        rom[278][13] = -8'd8;
        rom[278][14] = 8'd9;
        rom[278][15] = 8'd26;
        rom[278][16] = -8'd6;
        rom[278][17] = -8'd47;
        rom[278][18] = 8'd33;
        rom[278][19] = 8'd18;
        rom[278][20] = 8'd24;
        rom[278][21] = 8'd12;
        rom[278][22] = -8'd4;
        rom[278][23] = -8'd39;
        rom[278][24] = -8'd18;
        rom[278][25] = -8'd53;
        rom[278][26] = -8'd7;
        rom[278][27] = 8'd15;
        rom[278][28] = 8'd10;
        rom[278][29] = -8'd8;
        rom[278][30] = 8'd21;
        rom[278][31] = -8'd16;
        rom[279][0] = 8'd13;
        rom[279][1] = 8'd33;
        rom[279][2] = 8'd1;
        rom[279][3] = -8'd9;
        rom[279][4] = -8'd10;
        rom[279][5] = -8'd20;
        rom[279][6] = -8'd20;
        rom[279][7] = 8'd11;
        rom[279][8] = 8'd8;
        rom[279][9] = 8'd3;
        rom[279][10] = -8'd24;
        rom[279][11] = -8'd14;
        rom[279][12] = 8'd12;
        rom[279][13] = -8'd34;
        rom[279][14] = -8'd33;
        rom[279][15] = -8'd15;
        rom[279][16] = -8'd50;
        rom[279][17] = -8'd26;
        rom[279][18] = -8'd15;
        rom[279][19] = -8'd4;
        rom[279][20] = 8'd10;
        rom[279][21] = 8'd14;
        rom[279][22] = -8'd43;
        rom[279][23] = -8'd22;
        rom[279][24] = 8'd5;
        rom[279][25] = 8'd47;
        rom[279][26] = -8'd4;
        rom[279][27] = -8'd15;
        rom[279][28] = -8'd2;
        rom[279][29] = -8'd1;
        rom[279][30] = -8'd27;
        rom[279][31] = 8'd0;
        rom[280][0] = -8'd20;
        rom[280][1] = 8'd1;
        rom[280][2] = 8'd52;
        rom[280][3] = 8'd10;
        rom[280][4] = 8'd15;
        rom[280][5] = -8'd19;
        rom[280][6] = 8'd34;
        rom[280][7] = 8'd1;
        rom[280][8] = -8'd5;
        rom[280][9] = -8'd21;
        rom[280][10] = -8'd17;
        rom[280][11] = -8'd25;
        rom[280][12] = -8'd55;
        rom[280][13] = 8'd1;
        rom[280][14] = 8'd37;
        rom[280][15] = -8'd53;
        rom[280][16] = 8'd39;
        rom[280][17] = 8'd5;
        rom[280][18] = 8'd17;
        rom[280][19] = -8'd24;
        rom[280][20] = 8'd5;
        rom[280][21] = -8'd11;
        rom[280][22] = -8'd61;
        rom[280][23] = 8'd28;
        rom[280][24] = 8'd35;
        rom[280][25] = 8'd15;
        rom[280][26] = -8'd56;
        rom[280][27] = -8'd18;
        rom[280][28] = -8'd46;
        rom[280][29] = -8'd19;
        rom[280][30] = -8'd35;
        rom[280][31] = -8'd54;
        rom[281][0] = -8'd28;
        rom[281][1] = -8'd4;
        rom[281][2] = 8'd3;
        rom[281][3] = -8'd10;
        rom[281][4] = -8'd1;
        rom[281][5] = 8'd12;
        rom[281][6] = 8'd1;
        rom[281][7] = 8'd5;
        rom[281][8] = 8'd22;
        rom[281][9] = -8'd1;
        rom[281][10] = 8'd21;
        rom[281][11] = -8'd28;
        rom[281][12] = 8'd12;
        rom[281][13] = 8'd1;
        rom[281][14] = 8'd13;
        rom[281][15] = 8'd13;
        rom[281][16] = -8'd1;
        rom[281][17] = 8'd6;
        rom[281][18] = 8'd1;
        rom[281][19] = 8'd11;
        rom[281][20] = -8'd18;
        rom[281][21] = -8'd1;
        rom[281][22] = 8'd4;
        rom[281][23] = -8'd7;
        rom[281][24] = -8'd9;
        rom[281][25] = 8'd25;
        rom[281][26] = -8'd4;
        rom[281][27] = 8'd19;
        rom[281][28] = 8'd9;
        rom[281][29] = -8'd16;
        rom[281][30] = -8'd1;
        rom[281][31] = -8'd17;
        rom[282][0] = -8'd50;
        rom[282][1] = -8'd7;
        rom[282][2] = 8'd5;
        rom[282][3] = 8'd16;
        rom[282][4] = 8'd39;
        rom[282][5] = 8'd0;
        rom[282][6] = 8'd6;
        rom[282][7] = 8'd1;
        rom[282][8] = 8'd7;
        rom[282][9] = -8'd5;
        rom[282][10] = -8'd17;
        rom[282][11] = -8'd2;
        rom[282][12] = -8'd12;
        rom[282][13] = 8'd11;
        rom[282][14] = -8'd6;
        rom[282][15] = 8'd0;
        rom[282][16] = -8'd6;
        rom[282][17] = -8'd26;
        rom[282][18] = 8'd19;
        rom[282][19] = 8'd11;
        rom[282][20] = 8'd1;
        rom[282][21] = -8'd8;
        rom[282][22] = -8'd4;
        rom[282][23] = -8'd14;
        rom[282][24] = -8'd15;
        rom[282][25] = 8'd5;
        rom[282][26] = 8'd31;
        rom[282][27] = 8'd3;
        rom[282][28] = -8'd4;
        rom[282][29] = -8'd1;
        rom[282][30] = -8'd3;
        rom[282][31] = 8'd10;
        rom[283][0] = 8'd18;
        rom[283][1] = 8'd5;
        rom[283][2] = 8'd6;
        rom[283][3] = 8'd17;
        rom[283][4] = -8'd25;
        rom[283][5] = -8'd17;
        rom[283][6] = -8'd25;
        rom[283][7] = -8'd10;
        rom[283][8] = 8'd8;
        rom[283][9] = -8'd4;
        rom[283][10] = 8'd11;
        rom[283][11] = 8'd14;
        rom[283][12] = -8'd34;
        rom[283][13] = 8'd15;
        rom[283][14] = 8'd11;
        rom[283][15] = 8'd6;
        rom[283][16] = 8'd17;
        rom[283][17] = 8'd10;
        rom[283][18] = 8'd35;
        rom[283][19] = 8'd4;
        rom[283][20] = 8'd23;
        rom[283][21] = -8'd5;
        rom[283][22] = 8'd3;
        rom[283][23] = -8'd22;
        rom[283][24] = -8'd15;
        rom[283][25] = 8'd23;
        rom[283][26] = 8'd28;
        rom[283][27] = 8'd3;
        rom[283][28] = -8'd32;
        rom[283][29] = -8'd11;
        rom[283][30] = 8'd11;
        rom[283][31] = 8'd0;
        rom[284][0] = 8'd4;
        rom[284][1] = -8'd9;
        rom[284][2] = -8'd18;
        rom[284][3] = 8'd18;
        rom[284][4] = 8'd7;
        rom[284][5] = 8'd15;
        rom[284][6] = 8'd12;
        rom[284][7] = -8'd13;
        rom[284][8] = -8'd18;
        rom[284][9] = -8'd4;
        rom[284][10] = -8'd19;
        rom[284][11] = 8'd11;
        rom[284][12] = -8'd30;
        rom[284][13] = 8'd8;
        rom[284][14] = 8'd3;
        rom[284][15] = 8'd17;
        rom[284][16] = 8'd14;
        rom[284][17] = -8'd5;
        rom[284][18] = 8'd13;
        rom[284][19] = -8'd18;
        rom[284][20] = -8'd3;
        rom[284][21] = -8'd16;
        rom[284][22] = -8'd6;
        rom[284][23] = 8'd47;
        rom[284][24] = -8'd1;
        rom[284][25] = 8'd21;
        rom[284][26] = 8'd1;
        rom[284][27] = 8'd5;
        rom[284][28] = 8'd17;
        rom[284][29] = -8'd10;
        rom[284][30] = 8'd27;
        rom[284][31] = -8'd18;
        rom[285][0] = -8'd30;
        rom[285][1] = 8'd23;
        rom[285][2] = -8'd7;
        rom[285][3] = -8'd7;
        rom[285][4] = -8'd18;
        rom[285][5] = -8'd27;
        rom[285][6] = 8'd55;
        rom[285][7] = 8'd6;
        rom[285][8] = -8'd2;
        rom[285][9] = -8'd19;
        rom[285][10] = 8'd11;
        rom[285][11] = -8'd43;
        rom[285][12] = -8'd45;
        rom[285][13] = 8'd5;
        rom[285][14] = -8'd10;
        rom[285][15] = -8'd16;
        rom[285][16] = 8'd4;
        rom[285][17] = -8'd2;
        rom[285][18] = 8'd9;
        rom[285][19] = -8'd14;
        rom[285][20] = 8'd18;
        rom[285][21] = -8'd10;
        rom[285][22] = -8'd13;
        rom[285][23] = -8'd6;
        rom[285][24] = 8'd12;
        rom[285][25] = 8'd17;
        rom[285][26] = 8'd0;
        rom[285][27] = -8'd11;
        rom[285][28] = 8'd23;
        rom[285][29] = -8'd3;
        rom[285][30] = 8'd41;
        rom[285][31] = 8'd7;
        rom[286][0] = -8'd1;
        rom[286][1] = -8'd11;
        rom[286][2] = -8'd12;
        rom[286][3] = -8'd40;
        rom[286][4] = 8'd59;
        rom[286][5] = 8'd8;
        rom[286][6] = -8'd16;
        rom[286][7] = -8'd38;
        rom[286][8] = -8'd13;
        rom[286][9] = -8'd5;
        rom[286][10] = -8'd24;
        rom[286][11] = 8'd4;
        rom[286][12] = -8'd9;
        rom[286][13] = 8'd19;
        rom[286][14] = -8'd24;
        rom[286][15] = -8'd2;
        rom[286][16] = 8'd61;
        rom[286][17] = 8'd30;
        rom[286][18] = 8'd7;
        rom[286][19] = -8'd7;
        rom[286][20] = -8'd35;
        rom[286][21] = -8'd25;
        rom[286][22] = 8'd9;
        rom[286][23] = 8'd3;
        rom[286][24] = 8'd30;
        rom[286][25] = 8'd23;
        rom[286][26] = -8'd1;
        rom[286][27] = -8'd42;
        rom[286][28] = 8'd30;
        rom[286][29] = 8'd14;
        rom[286][30] = 8'd2;
        rom[286][31] = 8'd21;
        rom[287][0] = 8'd26;
        rom[287][1] = -8'd26;
        rom[287][2] = 8'd53;
        rom[287][3] = -8'd37;
        rom[287][4] = -8'd15;
        rom[287][5] = 8'd2;
        rom[287][6] = -8'd65;
        rom[287][7] = -8'd4;
        rom[287][8] = -8'd30;
        rom[287][9] = -8'd10;
        rom[287][10] = -8'd26;
        rom[287][11] = -8'd3;
        rom[287][12] = 8'd14;
        rom[287][13] = -8'd49;
        rom[287][14] = 8'd12;
        rom[287][15] = 8'd0;
        rom[287][16] = -8'd72;
        rom[287][17] = -8'd2;
        rom[287][18] = 8'd16;
        rom[287][19] = -8'd9;
        rom[287][20] = -8'd17;
        rom[287][21] = -8'd29;
        rom[287][22] = -8'd11;
        rom[287][23] = 8'd43;
        rom[287][24] = -8'd7;
        rom[287][25] = 8'd9;
        rom[287][26] = -8'd7;
        rom[287][27] = 8'd15;
        rom[287][28] = -8'd19;
        rom[287][29] = -8'd10;
        rom[287][30] = 8'd4;
        rom[287][31] = -8'd9;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
