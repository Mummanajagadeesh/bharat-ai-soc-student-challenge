module rom_01_conv2d_1_kernel (
    input  wire [15:0] row,
    input  wire [15:0] col,
    output reg signed [7:0] data
);

    // Q1.7 fixed-point format (8 bits total)
    reg signed [7:0] rom [0:143][0:15];

    initial begin
        rom[0][0] = 8'd8;
        rom[0][1] = -8'd14;
        rom[0][2] = -8'd9;
        rom[0][3] = 8'd11;
        rom[0][4] = 8'd17;
        rom[0][5] = -8'd9;
        rom[0][6] = -8'd6;
        rom[0][7] = 8'd7;
        rom[0][8] = -8'd8;
        rom[0][9] = 8'd8;
        rom[0][10] = 8'd13;
        rom[0][11] = 8'd15;
        rom[0][12] = -8'd7;
        rom[0][13] = 8'd13;
        rom[0][14] = 8'd18;
        rom[0][15] = 8'd11;
        rom[1][0] = 8'd25;
        rom[1][1] = -8'd39;
        rom[1][2] = 8'd10;
        rom[1][3] = -8'd7;
        rom[1][4] = 8'd8;
        rom[1][5] = -8'd17;
        rom[1][6] = -8'd31;
        rom[1][7] = 8'd17;
        rom[1][8] = -8'd7;
        rom[1][9] = 8'd2;
        rom[1][10] = -8'd24;
        rom[1][11] = 8'd24;
        rom[1][12] = -8'd11;
        rom[1][13] = -8'd5;
        rom[1][14] = 8'd17;
        rom[1][15] = 8'd14;
        rom[2][0] = -8'd34;
        rom[2][1] = -8'd18;
        rom[2][2] = 8'd33;
        rom[2][3] = -8'd27;
        rom[2][4] = -8'd45;
        rom[2][5] = -8'd7;
        rom[2][6] = 8'd7;
        rom[2][7] = 8'd29;
        rom[2][8] = -8'd19;
        rom[2][9] = 8'd12;
        rom[2][10] = 8'd16;
        rom[2][11] = -8'd24;
        rom[2][12] = -8'd22;
        rom[2][13] = -8'd49;
        rom[2][14] = -8'd11;
        rom[2][15] = -8'd12;
        rom[3][0] = 8'd31;
        rom[3][1] = 8'd8;
        rom[3][2] = 8'd1;
        rom[3][3] = 8'd12;
        rom[3][4] = 8'd25;
        rom[3][5] = 8'd49;
        rom[3][6] = 8'd7;
        rom[3][7] = 8'd22;
        rom[3][8] = -8'd18;
        rom[3][9] = -8'd17;
        rom[3][10] = -8'd15;
        rom[3][11] = -8'd16;
        rom[3][12] = -8'd15;
        rom[3][13] = 8'd13;
        rom[3][14] = -8'd3;
        rom[3][15] = -8'd7;
        rom[4][0] = -8'd59;
        rom[4][1] = -8'd10;
        rom[4][2] = -8'd12;
        rom[4][3] = 8'd11;
        rom[4][4] = 8'd23;
        rom[4][5] = -8'd11;
        rom[4][6] = 8'd1;
        rom[4][7] = -8'd17;
        rom[4][8] = -8'd25;
        rom[4][9] = -8'd17;
        rom[4][10] = -8'd6;
        rom[4][11] = 8'd20;
        rom[4][12] = 8'd7;
        rom[4][13] = 8'd2;
        rom[4][14] = -8'd2;
        rom[4][15] = -8'd13;
        rom[5][0] = -8'd4;
        rom[5][1] = -8'd17;
        rom[5][2] = 8'd16;
        rom[5][3] = -8'd11;
        rom[5][4] = -8'd34;
        rom[5][5] = -8'd1;
        rom[5][6] = 8'd13;
        rom[5][7] = -8'd17;
        rom[5][8] = 8'd10;
        rom[5][9] = -8'd1;
        rom[5][10] = -8'd1;
        rom[5][11] = -8'd5;
        rom[5][12] = 8'd16;
        rom[5][13] = -8'd16;
        rom[5][14] = -8'd2;
        rom[5][15] = 8'd17;
        rom[6][0] = 8'd23;
        rom[6][1] = 8'd41;
        rom[6][2] = 8'd30;
        rom[6][3] = 8'd69;
        rom[6][4] = 8'd26;
        rom[6][5] = 8'd4;
        rom[6][6] = -8'd9;
        rom[6][7] = -8'd20;
        rom[6][8] = 8'd9;
        rom[6][9] = -8'd4;
        rom[6][10] = 8'd14;
        rom[6][11] = 8'd13;
        rom[6][12] = 8'd18;
        rom[6][13] = -8'd8;
        rom[6][14] = 8'd8;
        rom[6][15] = 8'd6;
        rom[7][0] = -8'd10;
        rom[7][1] = -8'd14;
        rom[7][2] = -8'd37;
        rom[7][3] = 8'd6;
        rom[7][4] = 8'd4;
        rom[7][5] = 8'd14;
        rom[7][6] = -8'd10;
        rom[7][7] = -8'd3;
        rom[7][8] = -8'd26;
        rom[7][9] = 8'd40;
        rom[7][10] = 8'd12;
        rom[7][11] = 8'd8;
        rom[7][12] = -8'd2;
        rom[7][13] = -8'd45;
        rom[7][14] = -8'd12;
        rom[7][15] = -8'd23;
        rom[8][0] = -8'd54;
        rom[8][1] = -8'd9;
        rom[8][2] = 8'd3;
        rom[8][3] = 8'd18;
        rom[8][4] = -8'd23;
        rom[8][5] = -8'd22;
        rom[8][6] = -8'd18;
        rom[8][7] = -8'd24;
        rom[8][8] = 8'd69;
        rom[8][9] = 8'd23;
        rom[8][10] = 8'd14;
        rom[8][11] = 8'd23;
        rom[8][12] = -8'd18;
        rom[8][13] = 8'd7;
        rom[8][14] = 8'd39;
        rom[8][15] = -8'd6;
        rom[9][0] = 8'd58;
        rom[9][1] = -8'd57;
        rom[9][2] = -8'd3;
        rom[9][3] = 8'd11;
        rom[9][4] = 8'd14;
        rom[9][5] = 8'd18;
        rom[9][6] = -8'd48;
        rom[9][7] = -8'd10;
        rom[9][8] = -8'd26;
        rom[9][9] = 8'd4;
        rom[9][10] = -8'd6;
        rom[9][11] = -8'd21;
        rom[9][12] = 8'd9;
        rom[9][13] = 8'd19;
        rom[9][14] = 8'd4;
        rom[9][15] = -8'd30;
        rom[10][0] = 8'd1;
        rom[10][1] = -8'd24;
        rom[10][2] = 8'd10;
        rom[10][3] = 8'd5;
        rom[10][4] = 8'd1;
        rom[10][5] = 8'd8;
        rom[10][6] = -8'd26;
        rom[10][7] = -8'd9;
        rom[10][8] = -8'd21;
        rom[10][9] = 8'd6;
        rom[10][10] = -8'd23;
        rom[10][11] = -8'd10;
        rom[10][12] = -8'd79;
        rom[10][13] = 8'd2;
        rom[10][14] = -8'd13;
        rom[10][15] = 8'd12;
        rom[11][0] = -8'd24;
        rom[11][1] = -8'd8;
        rom[11][2] = -8'd26;
        rom[11][3] = 8'd10;
        rom[11][4] = 8'd29;
        rom[11][5] = -8'd2;
        rom[11][6] = 8'd9;
        rom[11][7] = 8'd6;
        rom[11][8] = 8'd2;
        rom[11][9] = -8'd14;
        rom[11][10] = 8'd9;
        rom[11][11] = 8'd28;
        rom[11][12] = 8'd40;
        rom[11][13] = 8'd8;
        rom[11][14] = 8'd30;
        rom[11][15] = 8'd26;
        rom[12][0] = -8'd31;
        rom[12][1] = -8'd9;
        rom[12][2] = -8'd27;
        rom[12][3] = -8'd7;
        rom[12][4] = -8'd9;
        rom[12][5] = 8'd7;
        rom[12][6] = -8'd18;
        rom[12][7] = 8'd17;
        rom[12][8] = 8'd3;
        rom[12][9] = -8'd2;
        rom[12][10] = -8'd2;
        rom[12][11] = 8'd16;
        rom[12][12] = 8'd25;
        rom[12][13] = -8'd5;
        rom[12][14] = -8'd2;
        rom[12][15] = 8'd20;
        rom[13][0] = -8'd14;
        rom[13][1] = -8'd6;
        rom[13][2] = 8'd39;
        rom[13][3] = 8'd0;
        rom[13][4] = 8'd9;
        rom[13][5] = 8'd11;
        rom[13][6] = 8'd11;
        rom[13][7] = 8'd14;
        rom[13][8] = -8'd16;
        rom[13][9] = -8'd2;
        rom[13][10] = 8'd41;
        rom[13][11] = -8'd36;
        rom[13][12] = 8'd3;
        rom[13][13] = -8'd41;
        rom[13][14] = 8'd5;
        rom[13][15] = -8'd68;
        rom[14][0] = 8'd16;
        rom[14][1] = -8'd20;
        rom[14][2] = 8'd33;
        rom[14][3] = 8'd57;
        rom[14][4] = 8'd29;
        rom[14][5] = 8'd53;
        rom[14][6] = 8'd19;
        rom[14][7] = -8'd3;
        rom[14][8] = -8'd1;
        rom[14][9] = -8'd24;
        rom[14][10] = 8'd10;
        rom[14][11] = 8'd6;
        rom[14][12] = 8'd45;
        rom[14][13] = -8'd7;
        rom[14][14] = -8'd38;
        rom[14][15] = -8'd32;
        rom[15][0] = 8'd32;
        rom[15][1] = 8'd71;
        rom[15][2] = 8'd4;
        rom[15][3] = 8'd23;
        rom[15][4] = 8'd6;
        rom[15][5] = -8'd11;
        rom[15][6] = -8'd6;
        rom[15][7] = -8'd23;
        rom[15][8] = -8'd22;
        rom[15][9] = -8'd26;
        rom[15][10] = -8'd5;
        rom[15][11] = -8'd51;
        rom[15][12] = -8'd19;
        rom[15][13] = 8'd11;
        rom[15][14] = 8'd49;
        rom[15][15] = -8'd23;
        rom[16][0] = 8'd2;
        rom[16][1] = -8'd18;
        rom[16][2] = -8'd22;
        rom[16][3] = 8'd3;
        rom[16][4] = -8'd17;
        rom[16][5] = -8'd3;
        rom[16][6] = -8'd8;
        rom[16][7] = 8'd2;
        rom[16][8] = -8'd6;
        rom[16][9] = -8'd3;
        rom[16][10] = 8'd17;
        rom[16][11] = 8'd6;
        rom[16][12] = 8'd15;
        rom[16][13] = 8'd16;
        rom[16][14] = 8'd14;
        rom[16][15] = -8'd2;
        rom[17][0] = 8'd16;
        rom[17][1] = 8'd1;
        rom[17][2] = 8'd20;
        rom[17][3] = -8'd16;
        rom[17][4] = 8'd8;
        rom[17][5] = 8'd5;
        rom[17][6] = -8'd25;
        rom[17][7] = 8'd4;
        rom[17][8] = -8'd18;
        rom[17][9] = 8'd15;
        rom[17][10] = 8'd3;
        rom[17][11] = -8'd47;
        rom[17][12] = -8'd46;
        rom[17][13] = 8'd26;
        rom[17][14] = -8'd29;
        rom[17][15] = -8'd12;
        rom[18][0] = -8'd11;
        rom[18][1] = -8'd44;
        rom[18][2] = 8'd0;
        rom[18][3] = -8'd16;
        rom[18][4] = -8'd5;
        rom[18][5] = -8'd3;
        rom[18][6] = -8'd7;
        rom[18][7] = -8'd26;
        rom[18][8] = 8'd7;
        rom[18][9] = -8'd20;
        rom[18][10] = -8'd16;
        rom[18][11] = -8'd45;
        rom[18][12] = 8'd7;
        rom[18][13] = -8'd8;
        rom[18][14] = -8'd19;
        rom[18][15] = 8'd5;
        rom[19][0] = 8'd22;
        rom[19][1] = -8'd1;
        rom[19][2] = -8'd28;
        rom[19][3] = 8'd8;
        rom[19][4] = 8'd53;
        rom[19][5] = -8'd56;
        rom[19][6] = -8'd21;
        rom[19][7] = 8'd1;
        rom[19][8] = 8'd21;
        rom[19][9] = -8'd72;
        rom[19][10] = -8'd36;
        rom[19][11] = 8'd38;
        rom[19][12] = 8'd14;
        rom[19][13] = -8'd1;
        rom[19][14] = 8'd57;
        rom[19][15] = -8'd3;
        rom[20][0] = 8'd1;
        rom[20][1] = 8'd15;
        rom[20][2] = -8'd51;
        rom[20][3] = 8'd26;
        rom[20][4] = 8'd20;
        rom[20][5] = 8'd5;
        rom[20][6] = 8'd3;
        rom[20][7] = 8'd1;
        rom[20][8] = -8'd29;
        rom[20][9] = 8'd36;
        rom[20][10] = -8'd48;
        rom[20][11] = 8'd20;
        rom[20][12] = -8'd4;
        rom[20][13] = 8'd11;
        rom[20][14] = 8'd22;
        rom[20][15] = 8'd30;
        rom[21][0] = 8'd7;
        rom[21][1] = 8'd10;
        rom[21][2] = -8'd9;
        rom[21][3] = 8'd12;
        rom[21][4] = -8'd27;
        rom[21][5] = 8'd28;
        rom[21][6] = -8'd1;
        rom[21][7] = -8'd23;
        rom[21][8] = 8'd10;
        rom[21][9] = 8'd23;
        rom[21][10] = 8'd10;
        rom[21][11] = -8'd22;
        rom[21][12] = 8'd10;
        rom[21][13] = 8'd5;
        rom[21][14] = -8'd30;
        rom[21][15] = -8'd27;
        rom[22][0] = 8'd11;
        rom[22][1] = 8'd21;
        rom[22][2] = -8'd7;
        rom[22][3] = 8'd18;
        rom[22][4] = 8'd22;
        rom[22][5] = -8'd17;
        rom[22][6] = 8'd11;
        rom[22][7] = -8'd14;
        rom[22][8] = -8'd2;
        rom[22][9] = -8'd35;
        rom[22][10] = 8'd14;
        rom[22][11] = -8'd1;
        rom[22][12] = 8'd12;
        rom[22][13] = -8'd12;
        rom[22][14] = 8'd23;
        rom[22][15] = -8'd19;
        rom[23][0] = 8'd9;
        rom[23][1] = 8'd6;
        rom[23][2] = -8'd24;
        rom[23][3] = -8'd3;
        rom[23][4] = -8'd2;
        rom[23][5] = -8'd1;
        rom[23][6] = 8'd1;
        rom[23][7] = 8'd19;
        rom[23][8] = -8'd33;
        rom[23][9] = 8'd22;
        rom[23][10] = 8'd10;
        rom[23][11] = -8'd11;
        rom[23][12] = -8'd21;
        rom[23][13] = -8'd21;
        rom[23][14] = 8'd4;
        rom[23][15] = -8'd1;
        rom[24][0] = -8'd36;
        rom[24][1] = -8'd5;
        rom[24][2] = 8'd37;
        rom[24][3] = 8'd14;
        rom[24][4] = 8'd5;
        rom[24][5] = 8'd5;
        rom[24][6] = 8'd10;
        rom[24][7] = 8'd6;
        rom[24][8] = 8'd2;
        rom[24][9] = 8'd23;
        rom[24][10] = 8'd55;
        rom[24][11] = -8'd42;
        rom[24][12] = 8'd12;
        rom[24][13] = 8'd3;
        rom[24][14] = -8'd13;
        rom[24][15] = -8'd37;
        rom[25][0] = 8'd64;
        rom[25][1] = -8'd10;
        rom[25][2] = -8'd7;
        rom[25][3] = -8'd4;
        rom[25][4] = 8'd28;
        rom[25][5] = -8'd20;
        rom[25][6] = -8'd42;
        rom[25][7] = -8'd2;
        rom[25][8] = -8'd42;
        rom[25][9] = -8'd16;
        rom[25][10] = -8'd23;
        rom[25][11] = 8'd20;
        rom[25][12] = -8'd4;
        rom[25][13] = 8'd12;
        rom[25][14] = -8'd6;
        rom[25][15] = -8'd8;
        rom[26][0] = 8'd20;
        rom[26][1] = 8'd13;
        rom[26][2] = 8'd3;
        rom[26][3] = -8'd1;
        rom[26][4] = -8'd7;
        rom[26][5] = -8'd26;
        rom[26][6] = -8'd42;
        rom[26][7] = 8'd5;
        rom[26][8] = -8'd15;
        rom[26][9] = -8'd15;
        rom[26][10] = 8'd17;
        rom[26][11] = -8'd16;
        rom[26][12] = 8'd6;
        rom[26][13] = -8'd27;
        rom[26][14] = -8'd23;
        rom[26][15] = -8'd15;
        rom[27][0] = -8'd17;
        rom[27][1] = 8'd24;
        rom[27][2] = 8'd19;
        rom[27][3] = 8'd13;
        rom[27][4] = 8'd52;
        rom[27][5] = -8'd15;
        rom[27][6] = 8'd5;
        rom[27][7] = -8'd30;
        rom[27][8] = 8'd11;
        rom[27][9] = -8'd40;
        rom[27][10] = -8'd31;
        rom[27][11] = 8'd22;
        rom[27][12] = 8'd64;
        rom[27][13] = -8'd6;
        rom[27][14] = -8'd47;
        rom[27][15] = 8'd6;
        rom[28][0] = -8'd27;
        rom[28][1] = -8'd28;
        rom[28][2] = 8'd48;
        rom[28][3] = 8'd2;
        rom[28][4] = -8'd10;
        rom[28][5] = -8'd43;
        rom[28][6] = 8'd0;
        rom[28][7] = -8'd22;
        rom[28][8] = 8'd20;
        rom[28][9] = -8'd22;
        rom[28][10] = 8'd32;
        rom[28][11] = 8'd10;
        rom[28][12] = 8'd1;
        rom[28][13] = 8'd27;
        rom[28][14] = 8'd22;
        rom[28][15] = -8'd18;
        rom[29][0] = -8'd16;
        rom[29][1] = 8'd23;
        rom[29][2] = -8'd3;
        rom[29][3] = 8'd6;
        rom[29][4] = 8'd1;
        rom[29][5] = -8'd19;
        rom[29][6] = 8'd10;
        rom[29][7] = 8'd20;
        rom[29][8] = 8'd8;
        rom[29][9] = -8'd14;
        rom[29][10] = -8'd3;
        rom[29][11] = 8'd12;
        rom[29][12] = -8'd3;
        rom[29][13] = -8'd12;
        rom[29][14] = -8'd56;
        rom[29][15] = 8'd16;
        rom[30][0] = -8'd15;
        rom[30][1] = -8'd37;
        rom[30][2] = -8'd38;
        rom[30][3] = 8'd38;
        rom[30][4] = 8'd23;
        rom[30][5] = -8'd37;
        rom[30][6] = 8'd18;
        rom[30][7] = 8'd26;
        rom[30][8] = 8'd8;
        rom[30][9] = -8'd39;
        rom[30][10] = 8'd29;
        rom[30][11] = 8'd54;
        rom[30][12] = 8'd51;
        rom[30][13] = -8'd15;
        rom[30][14] = -8'd1;
        rom[30][15] = 8'd34;
        rom[31][0] = 8'd34;
        rom[31][1] = 8'd83;
        rom[31][2] = -8'd9;
        rom[31][3] = 8'd10;
        rom[31][4] = -8'd6;
        rom[31][5] = -8'd42;
        rom[31][6] = -8'd20;
        rom[31][7] = 8'd4;
        rom[31][8] = -8'd44;
        rom[31][9] = -8'd10;
        rom[31][10] = -8'd13;
        rom[31][11] = -8'd7;
        rom[31][12] = 8'd13;
        rom[31][13] = 8'd2;
        rom[31][14] = -8'd21;
        rom[31][15] = -8'd17;
        rom[32][0] = -8'd1;
        rom[32][1] = 8'd11;
        rom[32][2] = 8'd13;
        rom[32][3] = 8'd4;
        rom[32][4] = 8'd2;
        rom[32][5] = 8'd6;
        rom[32][6] = -8'd19;
        rom[32][7] = 8'd16;
        rom[32][8] = 8'd19;
        rom[32][9] = -8'd20;
        rom[32][10] = -8'd11;
        rom[32][11] = 8'd19;
        rom[32][12] = 8'd6;
        rom[32][13] = -8'd8;
        rom[32][14] = 8'd9;
        rom[32][15] = -8'd8;
        rom[33][0] = 8'd39;
        rom[33][1] = 8'd16;
        rom[33][2] = 8'd0;
        rom[33][3] = 8'd11;
        rom[33][4] = 8'd19;
        rom[33][5] = 8'd8;
        rom[33][6] = -8'd44;
        rom[33][7] = 8'd11;
        rom[33][8] = -8'd13;
        rom[33][9] = 8'd10;
        rom[33][10] = -8'd1;
        rom[33][11] = 8'd18;
        rom[33][12] = -8'd27;
        rom[33][13] = 8'd8;
        rom[33][14] = 8'd9;
        rom[33][15] = 8'd0;
        rom[34][0] = -8'd15;
        rom[34][1] = -8'd100;
        rom[34][2] = -8'd15;
        rom[34][3] = 8'd15;
        rom[34][4] = -8'd7;
        rom[34][5] = 8'd16;
        rom[34][6] = 8'd5;
        rom[34][7] = -8'd16;
        rom[34][8] = 8'd5;
        rom[34][9] = 8'd36;
        rom[34][10] = -8'd16;
        rom[34][11] = -8'd30;
        rom[34][12] = 8'd7;
        rom[34][13] = 8'd11;
        rom[34][14] = -8'd30;
        rom[34][15] = 8'd37;
        rom[35][0] = -8'd1;
        rom[35][1] = 8'd0;
        rom[35][2] = 8'd46;
        rom[35][3] = 8'd15;
        rom[35][4] = 8'd42;
        rom[35][5] = 8'd1;
        rom[35][6] = 8'd18;
        rom[35][7] = -8'd24;
        rom[35][8] = 8'd37;
        rom[35][9] = 8'd1;
        rom[35][10] = 8'd9;
        rom[35][11] = -8'd54;
        rom[35][12] = 8'd47;
        rom[35][13] = 8'd8;
        rom[35][14] = -8'd10;
        rom[35][15] = -8'd9;
        rom[36][0] = 8'd6;
        rom[36][1] = 8'd4;
        rom[36][2] = 8'd13;
        rom[36][3] = 8'd35;
        rom[36][4] = 8'd20;
        rom[36][5] = -8'd3;
        rom[36][6] = 8'd13;
        rom[36][7] = 8'd32;
        rom[36][8] = -8'd31;
        rom[36][9] = -8'd30;
        rom[36][10] = -8'd2;
        rom[36][11] = -8'd11;
        rom[36][12] = -8'd3;
        rom[36][13] = -8'd25;
        rom[36][14] = -8'd17;
        rom[36][15] = -8'd1;
        rom[37][0] = 8'd23;
        rom[37][1] = 8'd19;
        rom[37][2] = -8'd9;
        rom[37][3] = 8'd4;
        rom[37][4] = -8'd34;
        rom[37][5] = -8'd11;
        rom[37][6] = 8'd6;
        rom[37][7] = -8'd3;
        rom[37][8] = -8'd5;
        rom[37][9] = 8'd7;
        rom[37][10] = 8'd5;
        rom[37][11] = 8'd27;
        rom[37][12] = 8'd18;
        rom[37][13] = -8'd19;
        rom[37][14] = -8'd18;
        rom[37][15] = 8'd9;
        rom[38][0] = 8'd17;
        rom[38][1] = -8'd37;
        rom[38][2] = 8'd1;
        rom[38][3] = -8'd10;
        rom[38][4] = 8'd46;
        rom[38][5] = 8'd13;
        rom[38][6] = 8'd6;
        rom[38][7] = -8'd27;
        rom[38][8] = 8'd19;
        rom[38][9] = 8'd13;
        rom[38][10] = -8'd17;
        rom[38][11] = -8'd27;
        rom[38][12] = 8'd10;
        rom[38][13] = 8'd13;
        rom[38][14] = 8'd32;
        rom[38][15] = 8'd2;
        rom[39][0] = -8'd11;
        rom[39][1] = 8'd14;
        rom[39][2] = 8'd26;
        rom[39][3] = -8'd21;
        rom[39][4] = -8'd28;
        rom[39][5] = -8'd34;
        rom[39][6] = 8'd3;
        rom[39][7] = 8'd14;
        rom[39][8] = -8'd4;
        rom[39][9] = 8'd1;
        rom[39][10] = 8'd10;
        rom[39][11] = -8'd17;
        rom[39][12] = 8'd0;
        rom[39][13] = -8'd12;
        rom[39][14] = 8'd35;
        rom[39][15] = 8'd36;
        rom[40][0] = 8'd3;
        rom[40][1] = -8'd6;
        rom[40][2] = -8'd31;
        rom[40][3] = 8'd22;
        rom[40][4] = -8'd12;
        rom[40][5] = -8'd1;
        rom[40][6] = 8'd26;
        rom[40][7] = 8'd29;
        rom[40][8] = -8'd27;
        rom[40][9] = -8'd41;
        rom[40][10] = -8'd40;
        rom[40][11] = 8'd17;
        rom[40][12] = 8'd5;
        rom[40][13] = -8'd33;
        rom[40][14] = 8'd33;
        rom[40][15] = 8'd30;
        rom[41][0] = 8'd4;
        rom[41][1] = -8'd48;
        rom[41][2] = -8'd7;
        rom[41][3] = -8'd55;
        rom[41][4] = 8'd15;
        rom[41][5] = -8'd49;
        rom[41][6] = -8'd4;
        rom[41][7] = -8'd21;
        rom[41][8] = -8'd22;
        rom[41][9] = -8'd37;
        rom[41][10] = -8'd28;
        rom[41][11] = -8'd14;
        rom[41][12] = 8'd45;
        rom[41][13] = 8'd49;
        rom[41][14] = -8'd3;
        rom[41][15] = 8'd7;
        rom[42][0] = -8'd18;
        rom[42][1] = 8'd43;
        rom[42][2] = -8'd32;
        rom[42][3] = -8'd12;
        rom[42][4] = 8'd7;
        rom[42][5] = 8'd7;
        rom[42][6] = -8'd19;
        rom[42][7] = -8'd4;
        rom[42][8] = -8'd7;
        rom[42][9] = -8'd27;
        rom[42][10] = -8'd15;
        rom[42][11] = 8'd7;
        rom[42][12] = 8'd22;
        rom[42][13] = 8'd22;
        rom[42][14] = 8'd2;
        rom[42][15] = -8'd8;
        rom[43][0] = -8'd5;
        rom[43][1] = 8'd7;
        rom[43][2] = -8'd6;
        rom[43][3] = 8'd30;
        rom[43][4] = 8'd44;
        rom[43][5] = -8'd6;
        rom[43][6] = -8'd1;
        rom[43][7] = -8'd46;
        rom[43][8] = -8'd6;
        rom[43][9] = -8'd24;
        rom[43][10] = 8'd2;
        rom[43][11] = -8'd23;
        rom[43][12] = 8'd21;
        rom[43][13] = 8'd8;
        rom[43][14] = -8'd71;
        rom[43][15] = -8'd25;
        rom[44][0] = -8'd20;
        rom[44][1] = -8'd11;
        rom[44][2] = -8'd14;
        rom[44][3] = 8'd28;
        rom[44][4] = -8'd12;
        rom[44][5] = 8'd2;
        rom[44][6] = 8'd9;
        rom[44][7] = -8'd52;
        rom[44][8] = 8'd29;
        rom[44][9] = 8'd9;
        rom[44][10] = 8'd16;
        rom[44][11] = -8'd29;
        rom[44][12] = 8'd7;
        rom[44][13] = 8'd39;
        rom[44][14] = 8'd4;
        rom[44][15] = -8'd21;
        rom[45][0] = -8'd29;
        rom[45][1] = -8'd16;
        rom[45][2] = -8'd28;
        rom[45][3] = 8'd6;
        rom[45][4] = 8'd5;
        rom[45][5] = -8'd4;
        rom[45][6] = 8'd16;
        rom[45][7] = 8'd13;
        rom[45][8] = 8'd8;
        rom[45][9] = -8'd13;
        rom[45][10] = -8'd41;
        rom[45][11] = 8'd3;
        rom[45][12] = 8'd27;
        rom[45][13] = -8'd32;
        rom[45][14] = -8'd13;
        rom[45][15] = 8'd33;
        rom[46][0] = -8'd24;
        rom[46][1] = -8'd20;
        rom[46][2] = -8'd16;
        rom[46][3] = 8'd49;
        rom[46][4] = 8'd36;
        rom[46][5] = 8'd9;
        rom[46][6] = 8'd49;
        rom[46][7] = -8'd9;
        rom[46][8] = 8'd18;
        rom[46][9] = -8'd49;
        rom[46][10] = -8'd31;
        rom[46][11] = -8'd20;
        rom[46][12] = 8'd8;
        rom[46][13] = -8'd14;
        rom[46][14] = -8'd34;
        rom[46][15] = 8'd21;
        rom[47][0] = 8'd6;
        rom[47][1] = 8'd1;
        rom[47][2] = 8'd16;
        rom[47][3] = -8'd1;
        rom[47][4] = -8'd17;
        rom[47][5] = -8'd10;
        rom[47][6] = 8'd4;
        rom[47][7] = -8'd9;
        rom[47][8] = -8'd20;
        rom[47][9] = -8'd29;
        rom[47][10] = 8'd30;
        rom[47][11] = -8'd6;
        rom[47][12] = -8'd13;
        rom[47][13] = 8'd6;
        rom[47][14] = 8'd5;
        rom[47][15] = -8'd6;
        rom[48][0] = 8'd8;
        rom[48][1] = -8'd1;
        rom[48][2] = -8'd6;
        rom[48][3] = 8'd16;
        rom[48][4] = 8'd6;
        rom[48][5] = 8'd8;
        rom[48][6] = 8'd2;
        rom[48][7] = -8'd8;
        rom[48][8] = -8'd15;
        rom[48][9] = -8'd8;
        rom[48][10] = 8'd7;
        rom[48][11] = -8'd1;
        rom[48][12] = -8'd2;
        rom[48][13] = 8'd11;
        rom[48][14] = 8'd3;
        rom[48][15] = 8'd11;
        rom[49][0] = 8'd18;
        rom[49][1] = -8'd38;
        rom[49][2] = -8'd2;
        rom[49][3] = 8'd16;
        rom[49][4] = 8'd2;
        rom[49][5] = -8'd31;
        rom[49][6] = 8'd29;
        rom[49][7] = -8'd25;
        rom[49][8] = 8'd11;
        rom[49][9] = 8'd5;
        rom[49][10] = 8'd16;
        rom[49][11] = 8'd0;
        rom[49][12] = -8'd41;
        rom[49][13] = -8'd21;
        rom[49][14] = 8'd18;
        rom[49][15] = 8'd20;
        rom[50][0] = -8'd12;
        rom[50][1] = 8'd42;
        rom[50][2] = -8'd16;
        rom[50][3] = 8'd5;
        rom[50][4] = -8'd21;
        rom[50][5] = 8'd11;
        rom[50][6] = 8'd22;
        rom[50][7] = -8'd7;
        rom[50][8] = 8'd43;
        rom[50][9] = -8'd17;
        rom[50][10] = 8'd17;
        rom[50][11] = -8'd10;
        rom[50][12] = 8'd17;
        rom[50][13] = -8'd22;
        rom[50][14] = -8'd16;
        rom[50][15] = -8'd19;
        rom[51][0] = -8'd43;
        rom[51][1] = -8'd3;
        rom[51][2] = 8'd31;
        rom[51][3] = 8'd28;
        rom[51][4] = -8'd31;
        rom[51][5] = 8'd46;
        rom[51][6] = -8'd2;
        rom[51][7] = 8'd27;
        rom[51][8] = 8'd51;
        rom[51][9] = -8'd45;
        rom[51][10] = 8'd47;
        rom[51][11] = -8'd4;
        rom[51][12] = -8'd8;
        rom[51][13] = 8'd0;
        rom[51][14] = -8'd34;
        rom[51][15] = -8'd35;
        rom[52][0] = 8'd26;
        rom[52][1] = -8'd5;
        rom[52][2] = 8'd18;
        rom[52][3] = -8'd38;
        rom[52][4] = -8'd11;
        rom[52][5] = 8'd23;
        rom[52][6] = 8'd18;
        rom[52][7] = -8'd11;
        rom[52][8] = -8'd15;
        rom[52][9] = 8'd16;
        rom[52][10] = 8'd16;
        rom[52][11] = -8'd23;
        rom[52][12] = 8'd7;
        rom[52][13] = -8'd35;
        rom[52][14] = -8'd16;
        rom[52][15] = -8'd52;
        rom[53][0] = -8'd11;
        rom[53][1] = -8'd1;
        rom[53][2] = -8'd12;
        rom[53][3] = 8'd11;
        rom[53][4] = 8'd17;
        rom[53][5] = -8'd19;
        rom[53][6] = 8'd1;
        rom[53][7] = -8'd62;
        rom[53][8] = -8'd14;
        rom[53][9] = 8'd2;
        rom[53][10] = -8'd18;
        rom[53][11] = -8'd6;
        rom[53][12] = -8'd4;
        rom[53][13] = 8'd10;
        rom[53][14] = 8'd3;
        rom[53][15] = 8'd9;
        rom[54][0] = -8'd30;
        rom[54][1] = 8'd43;
        rom[54][2] = -8'd15;
        rom[54][3] = 8'd43;
        rom[54][4] = -8'd11;
        rom[54][5] = -8'd6;
        rom[54][6] = -8'd1;
        rom[54][7] = 8'd13;
        rom[54][8] = 8'd29;
        rom[54][9] = -8'd14;
        rom[54][10] = -8'd26;
        rom[54][11] = 8'd28;
        rom[54][12] = -8'd4;
        rom[54][13] = 8'd7;
        rom[54][14] = 8'd1;
        rom[54][15] = 8'd30;
        rom[55][0] = 8'd22;
        rom[55][1] = 8'd3;
        rom[55][2] = -8'd26;
        rom[55][3] = -8'd6;
        rom[55][4] = -8'd21;
        rom[55][5] = 8'd36;
        rom[55][6] = -8'd16;
        rom[55][7] = 8'd24;
        rom[55][8] = 8'd19;
        rom[55][9] = 8'd14;
        rom[55][10] = -8'd10;
        rom[55][11] = 8'd8;
        rom[55][12] = -8'd34;
        rom[55][13] = -8'd48;
        rom[55][14] = 8'd12;
        rom[55][15] = 8'd12;
        rom[56][0] = 8'd1;
        rom[56][1] = -8'd3;
        rom[56][2] = -8'd27;
        rom[56][3] = 8'd12;
        rom[56][4] = 8'd37;
        rom[56][5] = 8'd0;
        rom[56][6] = -8'd19;
        rom[56][7] = -8'd18;
        rom[56][8] = -8'd59;
        rom[56][9] = 8'd10;
        rom[56][10] = -8'd73;
        rom[56][11] = 8'd33;
        rom[56][12] = -8'd15;
        rom[56][13] = 8'd6;
        rom[56][14] = 8'd37;
        rom[56][15] = 8'd38;
        rom[57][0] = 8'd9;
        rom[57][1] = 8'd5;
        rom[57][2] = -8'd7;
        rom[57][3] = 8'd5;
        rom[57][4] = 8'd7;
        rom[57][5] = 8'd33;
        rom[57][6] = 8'd9;
        rom[57][7] = 8'd24;
        rom[57][8] = 8'd0;
        rom[57][9] = 8'd14;
        rom[57][10] = -8'd8;
        rom[57][11] = -8'd18;
        rom[57][12] = -8'd13;
        rom[57][13] = 8'd24;
        rom[57][14] = 8'd8;
        rom[57][15] = 8'd3;
        rom[58][0] = 8'd38;
        rom[58][1] = -8'd25;
        rom[58][2] = -8'd1;
        rom[58][3] = 8'd35;
        rom[58][4] = -8'd7;
        rom[58][5] = 8'd20;
        rom[58][6] = 8'd23;
        rom[58][7] = 8'd16;
        rom[58][8] = -8'd15;
        rom[58][9] = -8'd20;
        rom[58][10] = -8'd19;
        rom[58][11] = 8'd1;
        rom[58][12] = -8'd38;
        rom[58][13] = -8'd12;
        rom[58][14] = -8'd10;
        rom[58][15] = 8'd16;
        rom[59][0] = 8'd22;
        rom[59][1] = 8'd28;
        rom[59][2] = -8'd14;
        rom[59][3] = -8'd34;
        rom[59][4] = -8'd29;
        rom[59][5] = -8'd8;
        rom[59][6] = 8'd30;
        rom[59][7] = 8'd15;
        rom[59][8] = 8'd31;
        rom[59][9] = 8'd0;
        rom[59][10] = 8'd18;
        rom[59][11] = -8'd15;
        rom[59][12] = 8'd8;
        rom[59][13] = 8'd19;
        rom[59][14] = 8'd27;
        rom[59][15] = -8'd2;
        rom[60][0] = -8'd7;
        rom[60][1] = -8'd8;
        rom[60][2] = -8'd36;
        rom[60][3] = 8'd0;
        rom[60][4] = -8'd3;
        rom[60][5] = -8'd12;
        rom[60][6] = 8'd3;
        rom[60][7] = -8'd3;
        rom[60][8] = -8'd14;
        rom[60][9] = 8'd9;
        rom[60][10] = -8'd22;
        rom[60][11] = 8'd28;
        rom[60][12] = 8'd0;
        rom[60][13] = 8'd16;
        rom[60][14] = -8'd5;
        rom[60][15] = 8'd32;
        rom[61][0] = 8'd8;
        rom[61][1] = 8'd19;
        rom[61][2] = 8'd9;
        rom[61][3] = 8'd3;
        rom[61][4] = -8'd12;
        rom[61][5] = 8'd25;
        rom[61][6] = -8'd11;
        rom[61][7] = 8'd28;
        rom[61][8] = -8'd1;
        rom[61][9] = -8'd36;
        rom[61][10] = -8'd11;
        rom[61][11] = -8'd8;
        rom[61][12] = -8'd20;
        rom[61][13] = -8'd40;
        rom[61][14] = 8'd22;
        rom[61][15] = -8'd46;
        rom[62][0] = 8'd0;
        rom[62][1] = 8'd18;
        rom[62][2] = 8'd28;
        rom[62][3] = -8'd27;
        rom[62][4] = 8'd18;
        rom[62][5] = 8'd24;
        rom[62][6] = -8'd41;
        rom[62][7] = 8'd31;
        rom[62][8] = -8'd11;
        rom[62][9] = -8'd37;
        rom[62][10] = -8'd5;
        rom[62][11] = -8'd20;
        rom[62][12] = 8'd48;
        rom[62][13] = 8'd9;
        rom[62][14] = 8'd8;
        rom[62][15] = -8'd19;
        rom[63][0] = 8'd31;
        rom[63][1] = 8'd64;
        rom[63][2] = 8'd1;
        rom[63][3] = -8'd24;
        rom[63][4] = -8'd20;
        rom[63][5] = -8'd17;
        rom[63][6] = 8'd19;
        rom[63][7] = 8'd3;
        rom[63][8] = -8'd23;
        rom[63][9] = -8'd26;
        rom[63][10] = 8'd7;
        rom[63][11] = -8'd35;
        rom[63][12] = 8'd7;
        rom[63][13] = -8'd3;
        rom[63][14] = 8'd43;
        rom[63][15] = -8'd19;
        rom[64][0] = -8'd15;
        rom[64][1] = -8'd15;
        rom[64][2] = 8'd2;
        rom[64][3] = 8'd0;
        rom[64][4] = 8'd0;
        rom[64][5] = 8'd22;
        rom[64][6] = 8'd10;
        rom[64][7] = 8'd9;
        rom[64][8] = -8'd6;
        rom[64][9] = 8'd1;
        rom[64][10] = 8'd9;
        rom[64][11] = -8'd6;
        rom[64][12] = 8'd5;
        rom[64][13] = 8'd3;
        rom[64][14] = -8'd5;
        rom[64][15] = 8'd9;
        rom[65][0] = 8'd35;
        rom[65][1] = -8'd22;
        rom[65][2] = -8'd2;
        rom[65][3] = 8'd8;
        rom[65][4] = -8'd22;
        rom[65][5] = 8'd41;
        rom[65][6] = 8'd2;
        rom[65][7] = -8'd3;
        rom[65][8] = 8'd20;
        rom[65][9] = -8'd11;
        rom[65][10] = -8'd14;
        rom[65][11] = -8'd65;
        rom[65][12] = -8'd45;
        rom[65][13] = 8'd22;
        rom[65][14] = -8'd7;
        rom[65][15] = -8'd16;
        rom[66][0] = -8'd28;
        rom[66][1] = 8'd32;
        rom[66][2] = -8'd1;
        rom[66][3] = 8'd1;
        rom[66][4] = -8'd18;
        rom[66][5] = -8'd17;
        rom[66][6] = 8'd28;
        rom[66][7] = -8'd60;
        rom[66][8] = 8'd21;
        rom[66][9] = 8'd21;
        rom[66][10] = 8'd12;
        rom[66][11] = -8'd12;
        rom[66][12] = 8'd15;
        rom[66][13] = 8'd17;
        rom[66][14] = 8'd0;
        rom[66][15] = -8'd26;
        rom[67][0] = -8'd28;
        rom[67][1] = -8'd10;
        rom[67][2] = -8'd46;
        rom[67][3] = 8'd25;
        rom[67][4] = -8'd40;
        rom[67][5] = -8'd86;
        rom[67][6] = 8'd22;
        rom[67][7] = -8'd40;
        rom[67][8] = 8'd49;
        rom[67][9] = 8'd5;
        rom[67][10] = 8'd11;
        rom[67][11] = 8'd37;
        rom[67][12] = 8'd17;
        rom[67][13] = 8'd11;
        rom[67][14] = 8'd21;
        rom[67][15] = 8'd31;
        rom[68][0] = 8'd3;
        rom[68][1] = -8'd7;
        rom[68][2] = -8'd21;
        rom[68][3] = 8'd6;
        rom[68][4] = 8'd15;
        rom[68][5] = -8'd24;
        rom[68][6] = 8'd4;
        rom[68][7] = 8'd33;
        rom[68][8] = 8'd23;
        rom[68][9] = -8'd38;
        rom[68][10] = 8'd19;
        rom[68][11] = -8'd5;
        rom[68][12] = 8'd16;
        rom[68][13] = 8'd9;
        rom[68][14] = -8'd8;
        rom[68][15] = 8'd24;
        rom[69][0] = 8'd20;
        rom[69][1] = 8'd12;
        rom[69][2] = -8'd7;
        rom[69][3] = 8'd21;
        rom[69][4] = 8'd22;
        rom[69][5] = 8'd31;
        rom[69][6] = -8'd15;
        rom[69][7] = 8'd8;
        rom[69][8] = -8'd22;
        rom[69][9] = 8'd13;
        rom[69][10] = -8'd17;
        rom[69][11] = -8'd28;
        rom[69][12] = 8'd3;
        rom[69][13] = -8'd8;
        rom[69][14] = 8'd4;
        rom[69][15] = -8'd9;
        rom[70][0] = -8'd13;
        rom[70][1] = 8'd28;
        rom[70][2] = -8'd15;
        rom[70][3] = 8'd20;
        rom[70][4] = -8'd21;
        rom[70][5] = 8'd5;
        rom[70][6] = -8'd19;
        rom[70][7] = -8'd29;
        rom[70][8] = 8'd9;
        rom[70][9] = 8'd20;
        rom[70][10] = 8'd13;
        rom[70][11] = -8'd6;
        rom[70][12] = 8'd8;
        rom[70][13] = -8'd28;
        rom[70][14] = 8'd30;
        rom[70][15] = -8'd60;
        rom[71][0] = 8'd1;
        rom[71][1] = 8'd22;
        rom[71][2] = -8'd46;
        rom[71][3] = -8'd23;
        rom[71][4] = -8'd27;
        rom[71][5] = -8'd40;
        rom[71][6] = -8'd23;
        rom[71][7] = 8'd3;
        rom[71][8] = 8'd16;
        rom[71][9] = 8'd8;
        rom[71][10] = 8'd8;
        rom[71][11] = 8'd20;
        rom[71][12] = -8'd39;
        rom[71][13] = -8'd31;
        rom[71][14] = 8'd2;
        rom[71][15] = -8'd18;
        rom[72][0] = 8'd25;
        rom[72][1] = 8'd18;
        rom[72][2] = 8'd44;
        rom[72][3] = 8'd5;
        rom[72][4] = 8'd35;
        rom[72][5] = 8'd25;
        rom[72][6] = -8'd77;
        rom[72][7] = 8'd24;
        rom[72][8] = -8'd56;
        rom[72][9] = -8'd1;
        rom[72][10] = 8'd3;
        rom[72][11] = -8'd51;
        rom[72][12] = -8'd1;
        rom[72][13] = 8'd5;
        rom[72][14] = -8'd33;
        rom[72][15] = -8'd63;
        rom[73][0] = -8'd46;
        rom[73][1] = 8'd14;
        rom[73][2] = -8'd5;
        rom[73][3] = 8'd1;
        rom[73][4] = 8'd37;
        rom[73][5] = -8'd29;
        rom[73][6] = -8'd32;
        rom[73][7] = -8'd16;
        rom[73][8] = 8'd3;
        rom[73][9] = -8'd41;
        rom[73][10] = -8'd24;
        rom[73][11] = 8'd3;
        rom[73][12] = 8'd19;
        rom[73][13] = 8'd4;
        rom[73][14] = -8'd19;
        rom[73][15] = -8'd21;
        rom[74][0] = 8'd0;
        rom[74][1] = -8'd17;
        rom[74][2] = -8'd8;
        rom[74][3] = 8'd25;
        rom[74][4] = 8'd6;
        rom[74][5] = -8'd29;
        rom[74][6] = -8'd2;
        rom[74][7] = -8'd19;
        rom[74][8] = 8'd14;
        rom[74][9] = -8'd10;
        rom[74][10] = 8'd14;
        rom[74][11] = -8'd27;
        rom[74][12] = 8'd5;
        rom[74][13] = -8'd41;
        rom[74][14] = -8'd2;
        rom[74][15] = 8'd9;
        rom[75][0] = 8'd5;
        rom[75][1] = 8'd49;
        rom[75][2] = 8'd12;
        rom[75][3] = -8'd56;
        rom[75][4] = -8'd2;
        rom[75][5] = -8'd25;
        rom[75][6] = 8'd32;
        rom[75][7] = -8'd27;
        rom[75][8] = 8'd6;
        rom[75][9] = 8'd17;
        rom[75][10] = 8'd0;
        rom[75][11] = 8'd15;
        rom[75][12] = 8'd34;
        rom[75][13] = -8'd3;
        rom[75][14] = -8'd16;
        rom[75][15] = 8'd19;
        rom[76][0] = 8'd9;
        rom[76][1] = 8'd4;
        rom[76][2] = -8'd3;
        rom[76][3] = -8'd21;
        rom[76][4] = -8'd5;
        rom[76][5] = -8'd15;
        rom[76][6] = -8'd14;
        rom[76][7] = -8'd87;
        rom[76][8] = -8'd22;
        rom[76][9] = 8'd31;
        rom[76][10] = -8'd45;
        rom[76][11] = -8'd1;
        rom[76][12] = 8'd7;
        rom[76][13] = 8'd35;
        rom[76][14] = 8'd33;
        rom[76][15] = 8'd21;
        rom[77][0] = -8'd26;
        rom[77][1] = 8'd49;
        rom[77][2] = 8'd39;
        rom[77][3] = 8'd3;
        rom[77][4] = -8'd10;
        rom[77][5] = -8'd6;
        rom[77][6] = 8'd10;
        rom[77][7] = 8'd16;
        rom[77][8] = 8'd20;
        rom[77][9] = -8'd8;
        rom[77][10] = 8'd32;
        rom[77][11] = 8'd9;
        rom[77][12] = -8'd3;
        rom[77][13] = -8'd29;
        rom[77][14] = -8'd50;
        rom[77][15] = -8'd24;
        rom[78][0] = -8'd19;
        rom[78][1] = 8'd40;
        rom[78][2] = 8'd10;
        rom[78][3] = -8'd30;
        rom[78][4] = 8'd31;
        rom[78][5] = -8'd70;
        rom[78][6] = -8'd65;
        rom[78][7] = -8'd8;
        rom[78][8] = 8'd4;
        rom[78][9] = -8'd31;
        rom[78][10] = 8'd31;
        rom[78][11] = 8'd7;
        rom[78][12] = 8'd42;
        rom[78][13] = 8'd19;
        rom[78][14] = 8'd24;
        rom[78][15] = 8'd1;
        rom[79][0] = 8'd49;
        rom[79][1] = 8'd89;
        rom[79][2] = -8'd12;
        rom[79][3] = -8'd1;
        rom[79][4] = -8'd1;
        rom[79][5] = -8'd11;
        rom[79][6] = -8'd15;
        rom[79][7] = -8'd18;
        rom[79][8] = -8'd25;
        rom[79][9] = 8'd10;
        rom[79][10] = -8'd8;
        rom[79][11] = -8'd15;
        rom[79][12] = 8'd3;
        rom[79][13] = -8'd3;
        rom[79][14] = -8'd29;
        rom[79][15] = -8'd4;
        rom[80][0] = -8'd12;
        rom[80][1] = -8'd6;
        rom[80][2] = -8'd11;
        rom[80][3] = -8'd10;
        rom[80][4] = 8'd16;
        rom[80][5] = -8'd6;
        rom[80][6] = 8'd1;
        rom[80][7] = 8'd4;
        rom[80][8] = -8'd4;
        rom[80][9] = -8'd11;
        rom[80][10] = 8'd0;
        rom[80][11] = 8'd10;
        rom[80][12] = 8'd9;
        rom[80][13] = 8'd9;
        rom[80][14] = 8'd10;
        rom[80][15] = -8'd18;
        rom[81][0] = 8'd32;
        rom[81][1] = 8'd19;
        rom[81][2] = -8'd11;
        rom[81][3] = 8'd9;
        rom[81][4] = 8'd0;
        rom[81][5] = -8'd15;
        rom[81][6] = 8'd5;
        rom[81][7] = 8'd4;
        rom[81][8] = 8'd27;
        rom[81][9] = -8'd29;
        rom[81][10] = -8'd13;
        rom[81][11] = 8'd26;
        rom[81][12] = -8'd1;
        rom[81][13] = -8'd4;
        rom[81][14] = 8'd15;
        rom[81][15] = -8'd14;
        rom[82][0] = 8'd50;
        rom[82][1] = -8'd5;
        rom[82][2] = -8'd3;
        rom[82][3] = -8'd21;
        rom[82][4] = -8'd32;
        rom[82][5] = 8'd8;
        rom[82][6] = 8'd19;
        rom[82][7] = -8'd24;
        rom[82][8] = 8'd13;
        rom[82][9] = -8'd7;
        rom[82][10] = 8'd15;
        rom[82][11] = 8'd20;
        rom[82][12] = -8'd15;
        rom[82][13] = -8'd28;
        rom[82][14] = -8'd12;
        rom[82][15] = 8'd19;
        rom[83][0] = -8'd37;
        rom[83][1] = -8'd8;
        rom[83][2] = 8'd31;
        rom[83][3] = -8'd14;
        rom[83][4] = -8'd39;
        rom[83][5] = 8'd39;
        rom[83][6] = 8'd18;
        rom[83][7] = -8'd12;
        rom[83][8] = -8'd11;
        rom[83][9] = 8'd11;
        rom[83][10] = -8'd22;
        rom[83][11] = -8'd65;
        rom[83][12] = 8'd9;
        rom[83][13] = 8'd14;
        rom[83][14] = -8'd2;
        rom[83][15] = 8'd6;
        rom[84][0] = 8'd27;
        rom[84][1] = 8'd8;
        rom[84][2] = 8'd17;
        rom[84][3] = 8'd23;
        rom[84][4] = -8'd7;
        rom[84][5] = -8'd3;
        rom[84][6] = -8'd25;
        rom[84][7] = -8'd5;
        rom[84][8] = 8'd18;
        rom[84][9] = -8'd38;
        rom[84][10] = -8'd6;
        rom[84][11] = 8'd0;
        rom[84][12] = 8'd9;
        rom[84][13] = 8'd1;
        rom[84][14] = -8'd35;
        rom[84][15] = -8'd10;
        rom[85][0] = -8'd3;
        rom[85][1] = 8'd35;
        rom[85][2] = -8'd6;
        rom[85][3] = 8'd30;
        rom[85][4] = 8'd15;
        rom[85][5] = -8'd27;
        rom[85][6] = 8'd0;
        rom[85][7] = 8'd19;
        rom[85][8] = -8'd20;
        rom[85][9] = -8'd27;
        rom[85][10] = 8'd21;
        rom[85][11] = 8'd34;
        rom[85][12] = 8'd6;
        rom[85][13] = 8'd9;
        rom[85][14] = -8'd14;
        rom[85][15] = -8'd18;
        rom[86][0] = -8'd4;
        rom[86][1] = 8'd11;
        rom[86][2] = -8'd22;
        rom[86][3] = -8'd30;
        rom[86][4] = -8'd27;
        rom[86][5] = 8'd13;
        rom[86][6] = 8'd9;
        rom[86][7] = 8'd3;
        rom[86][8] = 8'd20;
        rom[86][9] = 8'd39;
        rom[86][10] = 8'd6;
        rom[86][11] = -8'd11;
        rom[86][12] = -8'd19;
        rom[86][13] = -8'd14;
        rom[86][14] = 8'd31;
        rom[86][15] = -8'd6;
        rom[87][0] = 8'd7;
        rom[87][1] = 8'd30;
        rom[87][2] = 8'd18;
        rom[87][3] = -8'd24;
        rom[87][4] = -8'd13;
        rom[87][5] = -8'd10;
        rom[87][6] = -8'd34;
        rom[87][7] = -8'd13;
        rom[87][8] = 8'd24;
        rom[87][9] = 8'd36;
        rom[87][10] = 8'd18;
        rom[87][11] = -8'd12;
        rom[87][12] = 8'd15;
        rom[87][13] = -8'd25;
        rom[87][14] = 8'd18;
        rom[87][15] = 8'd11;
        rom[88][0] = -8'd5;
        rom[88][1] = 8'd7;
        rom[88][2] = -8'd7;
        rom[88][3] = -8'd32;
        rom[88][4] = 8'd21;
        rom[88][5] = -8'd29;
        rom[88][6] = -8'd29;
        rom[88][7] = 8'd9;
        rom[88][8] = 8'd12;
        rom[88][9] = 8'd1;
        rom[88][10] = 8'd59;
        rom[88][11] = 8'd25;
        rom[88][12] = 8'd18;
        rom[88][13] = -8'd4;
        rom[88][14] = -8'd11;
        rom[88][15] = 8'd9;
        rom[89][0] = -8'd14;
        rom[89][1] = 8'd9;
        rom[89][2] = -8'd1;
        rom[89][3] = -8'd6;
        rom[89][4] = 8'd31;
        rom[89][5] = -8'd5;
        rom[89][6] = -8'd4;
        rom[89][7] = 8'd16;
        rom[89][8] = -8'd11;
        rom[89][9] = -8'd27;
        rom[89][10] = -8'd39;
        rom[89][11] = -8'd24;
        rom[89][12] = 8'd18;
        rom[89][13] = 8'd22;
        rom[89][14] = -8'd7;
        rom[89][15] = 8'd8;
        rom[90][0] = -8'd4;
        rom[90][1] = 8'd16;
        rom[90][2] = 8'd10;
        rom[90][3] = 8'd6;
        rom[90][4] = 8'd11;
        rom[90][5] = 8'd26;
        rom[90][6] = -8'd26;
        rom[90][7] = 8'd4;
        rom[90][8] = 8'd6;
        rom[90][9] = 8'd20;
        rom[90][10] = 8'd7;
        rom[90][11] = 8'd5;
        rom[90][12] = 8'd39;
        rom[90][13] = -8'd2;
        rom[90][14] = -8'd19;
        rom[90][15] = -8'd25;
        rom[91][0] = -8'd6;
        rom[91][1] = 8'd45;
        rom[91][2] = 8'd5;
        rom[91][3] = -8'd29;
        rom[91][4] = -8'd8;
        rom[91][5] = 8'd17;
        rom[91][6] = 8'd12;
        rom[91][7] = -8'd7;
        rom[91][8] = -8'd9;
        rom[91][9] = 8'd0;
        rom[91][10] = -8'd17;
        rom[91][11] = 8'd0;
        rom[91][12] = -8'd12;
        rom[91][13] = 8'd1;
        rom[91][14] = -8'd36;
        rom[91][15] = -8'd22;
        rom[92][0] = -8'd24;
        rom[92][1] = 8'd7;
        rom[92][2] = 8'd14;
        rom[92][3] = -8'd5;
        rom[92][4] = -8'd6;
        rom[92][5] = 8'd44;
        rom[92][6] = -8'd13;
        rom[92][7] = -8'd21;
        rom[92][8] = -8'd37;
        rom[92][9] = 8'd33;
        rom[92][10] = -8'd9;
        rom[92][11] = -8'd16;
        rom[92][12] = -8'd17;
        rom[92][13] = 8'd10;
        rom[92][14] = -8'd5;
        rom[92][15] = -8'd20;
        rom[93][0] = 8'd32;
        rom[93][1] = 8'd5;
        rom[93][2] = -8'd39;
        rom[93][3] = -8'd11;
        rom[93][4] = -8'd19;
        rom[93][5] = -8'd5;
        rom[93][6] = 8'd3;
        rom[93][7] = -8'd4;
        rom[93][8] = 8'd2;
        rom[93][9] = 8'd32;
        rom[93][10] = 8'd19;
        rom[93][11] = 8'd3;
        rom[93][12] = 8'd14;
        rom[93][13] = -8'd24;
        rom[93][14] = 8'd24;
        rom[93][15] = 8'd36;
        rom[94][0] = -8'd39;
        rom[94][1] = 8'd41;
        rom[94][2] = -8'd28;
        rom[94][3] = -8'd10;
        rom[94][4] = 8'd14;
        rom[94][5] = 8'd42;
        rom[94][6] = -8'd9;
        rom[94][7] = -8'd33;
        rom[94][8] = -8'd15;
        rom[94][9] = 8'd24;
        rom[94][10] = 8'd7;
        rom[94][11] = -8'd58;
        rom[94][12] = -8'd6;
        rom[94][13] = 8'd11;
        rom[94][14] = -8'd12;
        rom[94][15] = 8'd30;
        rom[95][0] = 8'd20;
        rom[95][1] = 8'd0;
        rom[95][2] = -8'd5;
        rom[95][3] = -8'd10;
        rom[95][4] = 8'd27;
        rom[95][5] = -8'd20;
        rom[95][6] = 8'd16;
        rom[95][7] = -8'd20;
        rom[95][8] = 8'd0;
        rom[95][9] = -8'd4;
        rom[95][10] = 8'd19;
        rom[95][11] = -8'd3;
        rom[95][12] = -8'd2;
        rom[95][13] = -8'd3;
        rom[95][14] = 8'd5;
        rom[95][15] = 8'd4;
        rom[96][0] = -8'd5;
        rom[96][1] = -8'd18;
        rom[96][2] = -8'd3;
        rom[96][3] = -8'd11;
        rom[96][4] = -8'd13;
        rom[96][5] = 8'd6;
        rom[96][6] = -8'd8;
        rom[96][7] = 8'd14;
        rom[96][8] = -8'd9;
        rom[96][9] = 8'd7;
        rom[96][10] = 8'd12;
        rom[96][11] = -8'd7;
        rom[96][12] = -8'd3;
        rom[96][13] = -8'd10;
        rom[96][14] = 8'd10;
        rom[96][15] = 8'd14;
        rom[97][0] = 8'd21;
        rom[97][1] = -8'd63;
        rom[97][2] = 8'd6;
        rom[97][3] = 8'd15;
        rom[97][4] = -8'd10;
        rom[97][5] = 8'd5;
        rom[97][6] = -8'd12;
        rom[97][7] = 8'd23;
        rom[97][8] = 8'd11;
        rom[97][9] = 8'd7;
        rom[97][10] = -8'd2;
        rom[97][11] = 8'd20;
        rom[97][12] = -8'd44;
        rom[97][13] = -8'd15;
        rom[97][14] = 8'd4;
        rom[97][15] = 8'd4;
        rom[98][0] = -8'd26;
        rom[98][1] = 8'd12;
        rom[98][2] = 8'd11;
        rom[98][3] = 8'd8;
        rom[98][4] = 8'd29;
        rom[98][5] = -8'd10;
        rom[98][6] = 8'd5;
        rom[98][7] = -8'd9;
        rom[98][8] = -8'd32;
        rom[98][9] = 8'd33;
        rom[98][10] = 8'd29;
        rom[98][11] = 8'd22;
        rom[98][12] = 8'd16;
        rom[98][13] = -8'd2;
        rom[98][14] = -8'd56;
        rom[98][15] = -8'd4;
        rom[99][0] = -8'd20;
        rom[99][1] = 8'd1;
        rom[99][2] = 8'd8;
        rom[99][3] = 8'd18;
        rom[99][4] = 8'd12;
        rom[99][5] = -8'd15;
        rom[99][6] = -8'd31;
        rom[99][7] = -8'd18;
        rom[99][8] = -8'd35;
        rom[99][9] = 8'd35;
        rom[99][10] = -8'd35;
        rom[99][11] = -8'd12;
        rom[99][12] = -8'd1;
        rom[99][13] = 8'd2;
        rom[99][14] = -8'd37;
        rom[99][15] = -8'd38;
        rom[100][0] = 8'd25;
        rom[100][1] = -8'd8;
        rom[100][2] = 8'd21;
        rom[100][3] = -8'd35;
        rom[100][4] = -8'd35;
        rom[100][5] = 8'd37;
        rom[100][6] = -8'd7;
        rom[100][7] = 8'd23;
        rom[100][8] = 8'd11;
        rom[100][9] = 8'd0;
        rom[100][10] = -8'd22;
        rom[100][11] = 8'd11;
        rom[100][12] = -8'd30;
        rom[100][13] = -8'd44;
        rom[100][14] = 8'd21;
        rom[100][15] = -8'd22;
        rom[101][0] = -8'd7;
        rom[101][1] = -8'd17;
        rom[101][2] = 8'd29;
        rom[101][3] = 8'd24;
        rom[101][4] = 8'd28;
        rom[101][5] = 8'd13;
        rom[101][6] = -8'd17;
        rom[101][7] = -8'd14;
        rom[101][8] = -8'd8;
        rom[101][9] = 8'd0;
        rom[101][10] = 8'd23;
        rom[101][11] = 8'd4;
        rom[101][12] = -8'd33;
        rom[101][13] = -8'd15;
        rom[101][14] = 8'd18;
        rom[101][15] = 8'd20;
        rom[102][0] = -8'd16;
        rom[102][1] = -8'd21;
        rom[102][2] = -8'd23;
        rom[102][3] = 8'd12;
        rom[102][4] = 8'd2;
        rom[102][5] = -8'd10;
        rom[102][6] = -8'd9;
        rom[102][7] = 8'd8;
        rom[102][8] = -8'd42;
        rom[102][9] = -8'd2;
        rom[102][10] = 8'd6;
        rom[102][11] = 8'd6;
        rom[102][12] = 8'd12;
        rom[102][13] = 8'd21;
        rom[102][14] = -8'd45;
        rom[102][15] = 8'd91;
        rom[103][0] = -8'd2;
        rom[103][1] = -8'd37;
        rom[103][2] = 8'd16;
        rom[103][3] = -8'd15;
        rom[103][4] = 8'd0;
        rom[103][5] = -8'd1;
        rom[103][6] = 8'd29;
        rom[103][7] = 8'd20;
        rom[103][8] = -8'd12;
        rom[103][9] = 8'd0;
        rom[103][10] = 8'd18;
        rom[103][11] = -8'd6;
        rom[103][12] = -8'd22;
        rom[103][13] = -8'd5;
        rom[103][14] = -8'd13;
        rom[103][15] = 8'd12;
        rom[104][0] = 8'd34;
        rom[104][1] = -8'd37;
        rom[104][2] = -8'd29;
        rom[104][3] = -8'd2;
        rom[104][4] = -8'd26;
        rom[104][5] = 8'd26;
        rom[104][6] = 8'd32;
        rom[104][7] = 8'd15;
        rom[104][8] = 8'd26;
        rom[104][9] = -8'd46;
        rom[104][10] = 8'd48;
        rom[104][11] = -8'd13;
        rom[104][12] = 8'd0;
        rom[104][13] = 8'd6;
        rom[104][14] = 8'd4;
        rom[104][15] = 8'd34;
        rom[105][0] = -8'd73;
        rom[105][1] = -8'd15;
        rom[105][2] = -8'd6;
        rom[105][3] = -8'd40;
        rom[105][4] = -8'd36;
        rom[105][5] = 8'd17;
        rom[105][6] = 8'd17;
        rom[105][7] = 8'd16;
        rom[105][8] = -8'd1;
        rom[105][9] = 8'd53;
        rom[105][10] = 8'd25;
        rom[105][11] = -8'd6;
        rom[105][12] = 8'd36;
        rom[105][13] = -8'd3;
        rom[105][14] = 8'd13;
        rom[105][15] = -8'd8;
        rom[106][0] = 8'd1;
        rom[106][1] = -8'd38;
        rom[106][2] = 8'd16;
        rom[106][3] = -8'd49;
        rom[106][4] = 8'd12;
        rom[106][5] = -8'd14;
        rom[106][6] = 8'd20;
        rom[106][7] = 8'd11;
        rom[106][8] = -8'd6;
        rom[106][9] = 8'd1;
        rom[106][10] = -8'd28;
        rom[106][11] = 8'd15;
        rom[106][12] = 8'd14;
        rom[106][13] = 8'd15;
        rom[106][14] = 8'd21;
        rom[106][15] = 8'd16;
        rom[107][0] = 8'd31;
        rom[107][1] = 8'd2;
        rom[107][2] = -8'd6;
        rom[107][3] = 8'd4;
        rom[107][4] = -8'd48;
        rom[107][5] = -8'd4;
        rom[107][6] = -8'd21;
        rom[107][7] = 8'd26;
        rom[107][8] = -8'd21;
        rom[107][9] = 8'd29;
        rom[107][10] = -8'd13;
        rom[107][11] = -8'd9;
        rom[107][12] = -8'd3;
        rom[107][13] = 8'd1;
        rom[107][14] = 8'd56;
        rom[107][15] = 8'd6;
        rom[108][0] = 8'd21;
        rom[108][1] = -8'd59;
        rom[108][2] = 8'd23;
        rom[108][3] = 8'd22;
        rom[108][4] = 8'd1;
        rom[108][5] = 8'd0;
        rom[108][6] = 8'd19;
        rom[108][7] = -8'd45;
        rom[108][8] = -8'd6;
        rom[108][9] = 8'd25;
        rom[108][10] = 8'd26;
        rom[108][11] = -8'd2;
        rom[108][12] = -8'd2;
        rom[108][13] = 8'd20;
        rom[108][14] = -8'd42;
        rom[108][15] = -8'd2;
        rom[109][0] = -8'd4;
        rom[109][1] = -8'd7;
        rom[109][2] = -8'd6;
        rom[109][3] = 8'd3;
        rom[109][4] = 8'd6;
        rom[109][5] = 8'd0;
        rom[109][6] = -8'd33;
        rom[109][7] = 8'd19;
        rom[109][8] = -8'd23;
        rom[109][9] = -8'd28;
        rom[109][10] = -8'd14;
        rom[109][11] = -8'd9;
        rom[109][12] = -8'd14;
        rom[109][13] = 8'd4;
        rom[109][14] = 8'd40;
        rom[109][15] = 8'd5;
        rom[110][0] = -8'd1;
        rom[110][1] = -8'd31;
        rom[110][2] = 8'd6;
        rom[110][3] = -8'd60;
        rom[110][4] = -8'd42;
        rom[110][5] = -8'd17;
        rom[110][6] = 8'd17;
        rom[110][7] = 8'd0;
        rom[110][8] = -8'd9;
        rom[110][9] = 8'd3;
        rom[110][10] = 8'd3;
        rom[110][11] = -8'd43;
        rom[110][12] = 8'd8;
        rom[110][13] = -8'd7;
        rom[110][14] = -8'd27;
        rom[110][15] = -8'd10;
        rom[111][0] = 8'd19;
        rom[111][1] = -8'd5;
        rom[111][2] = 8'd15;
        rom[111][3] = -8'd18;
        rom[111][4] = 8'd2;
        rom[111][5] = -8'd21;
        rom[111][6] = 8'd6;
        rom[111][7] = 8'd21;
        rom[111][8] = -8'd25;
        rom[111][9] = -8'd8;
        rom[111][10] = 8'd22;
        rom[111][11] = -8'd52;
        rom[111][12] = 8'd9;
        rom[111][13] = -8'd20;
        rom[111][14] = 8'd26;
        rom[111][15] = -8'd5;
        rom[112][0] = 8'd4;
        rom[112][1] = 8'd3;
        rom[112][2] = -8'd17;
        rom[112][3] = -8'd3;
        rom[112][4] = 8'd19;
        rom[112][5] = -8'd8;
        rom[112][6] = 8'd14;
        rom[112][7] = 8'd15;
        rom[112][8] = -8'd8;
        rom[112][9] = 8'd0;
        rom[112][10] = -8'd16;
        rom[112][11] = -8'd9;
        rom[112][12] = -8'd10;
        rom[112][13] = 8'd2;
        rom[112][14] = -8'd16;
        rom[112][15] = 8'd9;
        rom[113][0] = 8'd6;
        rom[113][1] = -8'd45;
        rom[113][2] = -8'd16;
        rom[113][3] = 8'd0;
        rom[113][4] = -8'd3;
        rom[113][5] = 8'd17;
        rom[113][6] = 8'd32;
        rom[113][7] = -8'd10;
        rom[113][8] = -8'd16;
        rom[113][9] = -8'd8;
        rom[113][10] = 8'd12;
        rom[113][11] = -8'd27;
        rom[113][12] = 8'd2;
        rom[113][13] = 8'd27;
        rom[113][14] = -8'd24;
        rom[113][15] = 8'd28;
        rom[114][0] = -8'd12;
        rom[114][1] = 8'd29;
        rom[114][2] = 8'd9;
        rom[114][3] = 8'd5;
        rom[114][4] = 8'd44;
        rom[114][5] = 8'd15;
        rom[114][6] = -8'd14;
        rom[114][7] = 8'd0;
        rom[114][8] = -8'd40;
        rom[114][9] = -8'd11;
        rom[114][10] = -8'd16;
        rom[114][11] = 8'd26;
        rom[114][12] = -8'd1;
        rom[114][13] = 8'd6;
        rom[114][14] = -8'd38;
        rom[114][15] = -8'd35;
        rom[115][0] = -8'd19;
        rom[115][1] = -8'd2;
        rom[115][2] = -8'd25;
        rom[115][3] = -8'd13;
        rom[115][4] = 8'd6;
        rom[115][5] = -8'd11;
        rom[115][6] = -8'd46;
        rom[115][7] = -8'd11;
        rom[115][8] = -8'd80;
        rom[115][9] = 8'd43;
        rom[115][10] = 8'd27;
        rom[115][11] = 8'd40;
        rom[115][12] = 8'd3;
        rom[115][13] = 8'd9;
        rom[115][14] = 8'd2;
        rom[115][15] = -8'd22;
        rom[116][0] = -8'd1;
        rom[116][1] = 8'd15;
        rom[116][2] = 8'd21;
        rom[116][3] = -8'd42;
        rom[116][4] = -8'd34;
        rom[116][5] = -8'd56;
        rom[116][6] = -8'd25;
        rom[116][7] = 8'd3;
        rom[116][8] = 8'd40;
        rom[116][9] = 8'd15;
        rom[116][10] = 8'd14;
        rom[116][11] = 8'd4;
        rom[116][12] = -8'd22;
        rom[116][13] = 8'd8;
        rom[116][14] = 8'd6;
        rom[116][15] = 8'd4;
        rom[117][0] = 8'd12;
        rom[117][1] = 8'd11;
        rom[117][2] = -8'd16;
        rom[117][3] = 8'd43;
        rom[117][4] = -8'd1;
        rom[117][5] = 8'd1;
        rom[117][6] = 8'd11;
        rom[117][7] = 8'd11;
        rom[117][8] = 8'd17;
        rom[117][9] = -8'd18;
        rom[117][10] = -8'd1;
        rom[117][11] = -8'd31;
        rom[117][12] = -8'd4;
        rom[117][13] = 8'd7;
        rom[117][14] = 8'd7;
        rom[117][15] = 8'd13;
        rom[118][0] = 8'd1;
        rom[118][1] = 8'd5;
        rom[118][2] = -8'd31;
        rom[118][3] = -8'd18;
        rom[118][4] = 8'd17;
        rom[118][5] = -8'd3;
        rom[118][6] = -8'd20;
        rom[118][7] = 8'd18;
        rom[118][8] = -8'd24;
        rom[118][9] = 8'd21;
        rom[118][10] = -8'd46;
        rom[118][11] = 8'd20;
        rom[118][12] = 8'd7;
        rom[118][13] = 8'd9;
        rom[118][14] = -8'd20;
        rom[118][15] = -8'd31;
        rom[119][0] = 8'd2;
        rom[119][1] = 8'd10;
        rom[119][2] = -8'd65;
        rom[119][3] = 8'd13;
        rom[119][4] = 8'd0;
        rom[119][5] = -8'd22;
        rom[119][6] = 8'd7;
        rom[119][7] = -8'd38;
        rom[119][8] = 8'd13;
        rom[119][9] = 8'd17;
        rom[119][10] = -8'd42;
        rom[119][11] = 8'd9;
        rom[119][12] = -8'd6;
        rom[119][13] = 8'd1;
        rom[119][14] = -8'd22;
        rom[119][15] = -8'd17;
        rom[120][0] = 8'd16;
        rom[120][1] = -8'd16;
        rom[120][2] = -8'd21;
        rom[120][3] = -8'd20;
        rom[120][4] = -8'd30;
        rom[120][5] = 8'd4;
        rom[120][6] = 8'd39;
        rom[120][7] = 8'd20;
        rom[120][8] = 8'd36;
        rom[120][9] = -8'd52;
        rom[120][10] = -8'd64;
        rom[120][11] = -8'd30;
        rom[120][12] = 8'd20;
        rom[120][13] = 8'd15;
        rom[120][14] = 8'd12;
        rom[120][15] = 8'd3;
        rom[121][0] = -8'd40;
        rom[121][1] = 8'd9;
        rom[121][2] = -8'd19;
        rom[121][3] = -8'd13;
        rom[121][4] = -8'd31;
        rom[121][5] = -8'd2;
        rom[121][6] = 8'd24;
        rom[121][7] = -8'd10;
        rom[121][8] = 8'd3;
        rom[121][9] = 8'd39;
        rom[121][10] = 8'd41;
        rom[121][11] = 8'd10;
        rom[121][12] = 8'd13;
        rom[121][13] = 8'd1;
        rom[121][14] = 8'd21;
        rom[121][15] = -8'd13;
        rom[122][0] = 8'd10;
        rom[122][1] = 8'd8;
        rom[122][2] = -8'd43;
        rom[122][3] = -8'd26;
        rom[122][4] = 8'd3;
        rom[122][5] = -8'd3;
        rom[122][6] = 8'd48;
        rom[122][7] = -8'd35;
        rom[122][8] = 8'd15;
        rom[122][9] = 8'd50;
        rom[122][10] = -8'd27;
        rom[122][11] = -8'd2;
        rom[122][12] = 8'd23;
        rom[122][13] = -8'd29;
        rom[122][14] = 8'd19;
        rom[122][15] = 8'd37;
        rom[123][0] = 8'd24;
        rom[123][1] = 8'd11;
        rom[123][2] = -8'd5;
        rom[123][3] = -8'd15;
        rom[123][4] = -8'd32;
        rom[123][5] = 8'd7;
        rom[123][6] = -8'd1;
        rom[123][7] = -8'd23;
        rom[123][8] = 8'd6;
        rom[123][9] = 8'd40;
        rom[123][10] = 8'd7;
        rom[123][11] = 8'd8;
        rom[123][12] = -8'd11;
        rom[123][13] = 8'd0;
        rom[123][14] = 8'd12;
        rom[123][15] = 8'd15;
        rom[124][0] = 8'd21;
        rom[124][1] = -8'd40;
        rom[124][2] = -8'd17;
        rom[124][3] = -8'd4;
        rom[124][4] = -8'd6;
        rom[124][5] = -8'd13;
        rom[124][6] = -8'd1;
        rom[124][7] = -8'd18;
        rom[124][8] = 8'd12;
        rom[124][9] = 8'd5;
        rom[124][10] = 8'd3;
        rom[124][11] = 8'd11;
        rom[124][12] = -8'd28;
        rom[124][13] = 8'd12;
        rom[124][14] = 8'd14;
        rom[124][15] = 8'd40;
        rom[125][0] = -8'd20;
        rom[125][1] = 8'd15;
        rom[125][2] = 8'd31;
        rom[125][3] = -8'd5;
        rom[125][4] = 8'd1;
        rom[125][5] = -8'd11;
        rom[125][6] = -8'd17;
        rom[125][7] = -8'd1;
        rom[125][8] = -8'd7;
        rom[125][9] = 8'd11;
        rom[125][10] = -8'd21;
        rom[125][11] = -8'd5;
        rom[125][12] = 8'd4;
        rom[125][13] = -8'd6;
        rom[125][14] = -8'd16;
        rom[125][15] = -8'd43;
        rom[126][0] = 8'd29;
        rom[126][1] = 8'd17;
        rom[126][2] = 8'd21;
        rom[126][3] = -8'd92;
        rom[126][4] = -8'd43;
        rom[126][5] = -8'd25;
        rom[126][6] = -8'd49;
        rom[126][7] = -8'd11;
        rom[126][8] = -8'd10;
        rom[126][9] = 8'd19;
        rom[126][10] = -8'd25;
        rom[126][11] = 8'd22;
        rom[126][12] = -8'd23;
        rom[126][13] = 8'd19;
        rom[126][14] = -8'd25;
        rom[126][15] = -8'd19;
        rom[127][0] = 8'd44;
        rom[127][1] = 8'd61;
        rom[127][2] = -8'd17;
        rom[127][3] = -8'd1;
        rom[127][4] = -8'd11;
        rom[127][5] = -8'd23;
        rom[127][6] = -8'd10;
        rom[127][7] = -8'd21;
        rom[127][8] = -8'd12;
        rom[127][9] = 8'd0;
        rom[127][10] = 8'd10;
        rom[127][11] = 8'd3;
        rom[127][12] = -8'd10;
        rom[127][13] = 8'd19;
        rom[127][14] = -8'd14;
        rom[127][15] = 8'd17;
        rom[128][0] = -8'd8;
        rom[128][1] = -8'd7;
        rom[128][2] = -8'd17;
        rom[128][3] = 8'd20;
        rom[128][4] = -8'd12;
        rom[128][5] = -8'd14;
        rom[128][6] = -8'd10;
        rom[128][7] = 8'd10;
        rom[128][8] = -8'd21;
        rom[128][9] = 8'd7;
        rom[128][10] = -8'd12;
        rom[128][11] = -8'd9;
        rom[128][12] = -8'd15;
        rom[128][13] = -8'd5;
        rom[128][14] = -8'd8;
        rom[128][15] = 8'd1;
        rom[129][0] = 8'd6;
        rom[129][1] = 8'd0;
        rom[129][2] = 8'd7;
        rom[129][3] = -8'd1;
        rom[129][4] = 8'd2;
        rom[129][5] = -8'd17;
        rom[129][6] = 8'd29;
        rom[129][7] = 8'd9;
        rom[129][8] = -8'd29;
        rom[129][9] = -8'd9;
        rom[129][10] = 8'd6;
        rom[129][11] = 8'd28;
        rom[129][12] = 8'd13;
        rom[129][13] = 8'd16;
        rom[129][14] = -8'd7;
        rom[129][15] = -8'd18;
        rom[130][0] = -8'd30;
        rom[130][1] = -8'd9;
        rom[130][2] = 8'd7;
        rom[130][3] = 8'd4;
        rom[130][4] = 8'd13;
        rom[130][5] = -8'd23;
        rom[130][6] = -8'd50;
        rom[130][7] = 8'd6;
        rom[130][8] = -8'd32;
        rom[130][9] = -8'd2;
        rom[130][10] = -8'd18;
        rom[130][11] = 8'd5;
        rom[130][12] = -8'd23;
        rom[130][13] = -8'd37;
        rom[130][14] = -8'd40;
        rom[130][15] = 8'd8;
        rom[131][0] = -8'd25;
        rom[131][1] = 8'd2;
        rom[131][2] = -8'd15;
        rom[131][3] = -8'd28;
        rom[131][4] = -8'd8;
        rom[131][5] = 8'd41;
        rom[131][6] = -8'd7;
        rom[131][7] = 8'd7;
        rom[131][8] = -8'd49;
        rom[131][9] = -8'd21;
        rom[131][10] = 8'd20;
        rom[131][11] = -8'd32;
        rom[131][12] = 8'd3;
        rom[131][13] = -8'd8;
        rom[131][14] = 8'd0;
        rom[131][15] = 8'd34;
        rom[132][0] = -8'd1;
        rom[132][1] = -8'd6;
        rom[132][2] = 8'd4;
        rom[132][3] = 8'd24;
        rom[132][4] = -8'd5;
        rom[132][5] = 8'd28;
        rom[132][6] = -8'd17;
        rom[132][7] = -8'd27;
        rom[132][8] = -8'd5;
        rom[132][9] = 8'd41;
        rom[132][10] = 8'd16;
        rom[132][11] = 8'd6;
        rom[132][12] = -8'd20;
        rom[132][13] = 8'd30;
        rom[132][14] = 8'd8;
        rom[132][15] = 8'd22;
        rom[133][0] = -8'd1;
        rom[133][1] = 8'd19;
        rom[133][2] = 8'd4;
        rom[133][3] = 8'd43;
        rom[133][4] = 8'd0;
        rom[133][5] = -8'd8;
        rom[133][6] = -8'd25;
        rom[133][7] = 8'd42;
        rom[133][8] = 8'd9;
        rom[133][9] = -8'd1;
        rom[133][10] = -8'd14;
        rom[133][11] = 8'd10;
        rom[133][12] = 8'd2;
        rom[133][13] = -8'd25;
        rom[133][14] = -8'd12;
        rom[133][15] = -8'd5;
        rom[134][0] = -8'd3;
        rom[134][1] = -8'd8;
        rom[134][2] = -8'd53;
        rom[134][3] = -8'd59;
        rom[134][4] = -8'd6;
        rom[134][5] = 8'd1;
        rom[134][6] = -8'd30;
        rom[134][7] = 8'd32;
        rom[134][8] = -8'd18;
        rom[134][9] = -8'd12;
        rom[134][10] = 8'd29;
        rom[134][11] = -8'd12;
        rom[134][12] = -8'd17;
        rom[134][13] = 8'd25;
        rom[134][14] = 8'd4;
        rom[134][15] = -8'd57;
        rom[135][0] = 8'd27;
        rom[135][1] = 8'd22;
        rom[135][2] = 8'd8;
        rom[135][3] = 8'd14;
        rom[135][4] = 8'd20;
        rom[135][5] = 8'd36;
        rom[135][6] = -8'd6;
        rom[135][7] = 8'd8;
        rom[135][8] = -8'd23;
        rom[135][9] = -8'd4;
        rom[135][10] = -8'd6;
        rom[135][11] = -8'd10;
        rom[135][12] = 8'd13;
        rom[135][13] = -8'd16;
        rom[135][14] = 8'd12;
        rom[135][15] = -8'd11;
        rom[136][0] = 8'd7;
        rom[136][1] = 8'd22;
        rom[136][2] = 8'd39;
        rom[136][3] = -8'd13;
        rom[136][4] = -8'd12;
        rom[136][5] = -8'd16;
        rom[136][6] = -8'd27;
        rom[136][7] = -8'd17;
        rom[136][8] = 8'd20;
        rom[136][9] = 8'd50;
        rom[136][10] = -8'd12;
        rom[136][11] = 8'd5;
        rom[136][12] = 8'd19;
        rom[136][13] = -8'd12;
        rom[136][14] = -8'd8;
        rom[136][15] = -8'd17;
        rom[137][0] = 8'd28;
        rom[137][1] = 8'd7;
        rom[137][2] = 8'd8;
        rom[137][3] = -8'd9;
        rom[137][4] = -8'd25;
        rom[137][5] = 8'd9;
        rom[137][6] = 8'd24;
        rom[137][7] = 8'd18;
        rom[137][8] = 8'd24;
        rom[137][9] = 8'd11;
        rom[137][10] = -8'd16;
        rom[137][11] = 8'd6;
        rom[137][12] = -8'd12;
        rom[137][13] = -8'd18;
        rom[137][14] = 8'd17;
        rom[137][15] = 8'd5;
        rom[138][0] = -8'd18;
        rom[138][1] = 8'd13;
        rom[138][2] = 8'd14;
        rom[138][3] = 8'd12;
        rom[138][4] = 8'd7;
        rom[138][5] = 8'd10;
        rom[138][6] = 8'd33;
        rom[138][7] = 8'd3;
        rom[138][8] = -8'd4;
        rom[138][9] = 8'd2;
        rom[138][10] = -8'd27;
        rom[138][11] = -8'd2;
        rom[138][12] = 8'd33;
        rom[138][13] = 8'd13;
        rom[138][14] = 8'd26;
        rom[138][15] = -8'd21;
        rom[139][0] = -8'd1;
        rom[139][1] = 8'd24;
        rom[139][2] = 8'd26;
        rom[139][3] = -8'd26;
        rom[139][4] = -8'd22;
        rom[139][5] = 8'd24;
        rom[139][6] = 8'd4;
        rom[139][7] = 8'd10;
        rom[139][8] = -8'd30;
        rom[139][9] = 8'd35;
        rom[139][10] = 8'd11;
        rom[139][11] = 8'd11;
        rom[139][12] = -8'd35;
        rom[139][13] = -8'd3;
        rom[139][14] = -8'd3;
        rom[139][15] = 8'd20;
        rom[140][0] = 8'd7;
        rom[140][1] = -8'd45;
        rom[140][2] = -8'd6;
        rom[140][3] = 8'd1;
        rom[140][4] = 8'd0;
        rom[140][5] = 8'd23;
        rom[140][6] = -8'd3;
        rom[140][7] = -8'd7;
        rom[140][8] = 8'd22;
        rom[140][9] = -8'd12;
        rom[140][10] = -8'd17;
        rom[140][11] = -8'd11;
        rom[140][12] = -8'd15;
        rom[140][13] = 8'd21;
        rom[140][14] = -8'd8;
        rom[140][15] = -8'd26;
        rom[141][0] = 8'd23;
        rom[141][1] = -8'd5;
        rom[141][2] = 8'd19;
        rom[141][3] = 8'd5;
        rom[141][4] = 8'd17;
        rom[141][5] = 8'd0;
        rom[141][6] = -8'd11;
        rom[141][7] = 8'd16;
        rom[141][8] = -8'd4;
        rom[141][9] = 8'd9;
        rom[141][10] = 8'd4;
        rom[141][11] = 8'd17;
        rom[141][12] = -8'd26;
        rom[141][13] = -8'd48;
        rom[141][14] = -8'd11;
        rom[141][15] = 8'd24;
        rom[142][0] = 8'd37;
        rom[142][1] = 8'd6;
        rom[142][2] = 8'd2;
        rom[142][3] = -8'd26;
        rom[142][4] = -8'd42;
        rom[142][5] = 8'd36;
        rom[142][6] = -8'd31;
        rom[142][7] = -8'd12;
        rom[142][8] = -8'd9;
        rom[142][9] = 8'd22;
        rom[142][10] = -8'd1;
        rom[142][11] = -8'd29;
        rom[142][12] = -8'd59;
        rom[142][13] = -8'd16;
        rom[142][14] = -8'd49;
        rom[142][15] = -8'd17;
        rom[143][0] = 8'd9;
        rom[143][1] = 8'd7;
        rom[143][2] = 8'd5;
        rom[143][3] = -8'd23;
        rom[143][4] = -8'd7;
        rom[143][5] = 8'd7;
        rom[143][6] = 8'd0;
        rom[143][7] = 8'd23;
        rom[143][8] = -8'd7;
        rom[143][9] = -8'd17;
        rom[143][10] = -8'd4;
        rom[143][11] = 8'd2;
        rom[143][12] = -8'd14;
        rom[143][13] = -8'd8;
        rom[143][14] = -8'd4;
        rom[143][15] = 8'd15;
    end

    always @(*) begin
        data = rom[row][col];
    end

endmodule
